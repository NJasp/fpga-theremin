library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
-- TESTFILE | proof of concept,
-- this will be done by the C code eventually hopefully
-- write induvidual sinus values to play any sinus wave

entity testFile is
port (
  CLOCK_50, CLOCK_27 : in std_logic;
  KEY : in std_logic_vector(3 downto 0);
  AUD_ADCDAT : in std_logic;
  AUD_BCLK : inout std_logic;
  AUD_ADCLRCK : inout std_logic;
  AUD_DACLRCK : inout std_logic;
  I2C_SDAT : inout std_logic;
  AUD_XCK : out std_logic;
  AUD_DACDAT : out std_logic;
  I2C_SCLK : out std_logic;
  LEDR : out std_logic_vector(17 downto 0);
  SW : in std_logic_vector(17 downto 0)
);
end testFile;

architecture behaviour of testFile is
	component DE2_Audio_Example port (
	  sinVal : in signed(13 downto 0);
	  CLOCK_50, CLOCK_27 : in std_logic;
	  KEY : in std_logic_vector(3 downto 0);
	  AUD_ADCDAT : in std_logic;
	  AUD_BCLK : inout std_logic;
	  AUD_ADCLRCK : inout std_logic;
	  AUD_DACLRCK : inout std_logic;
	  I2C_SDAT : inout std_logic;
	  AUD_XCK : out std_logic;
	  AUD_DACDAT : out std_logic;
	  I2C_SCLK : out std_logic;
	  LEDR : out std_logic_vector(17 downto 0);
	  SW : in std_logic_vector(17 downto 0)
	);
	end component;
	
	signal delay_cnt, delay : signed(18 downto 0);
	signal acc : unsigned(8 downto 0);
	signal sinVal : signed(13 downto 0);
	
begin
	process(CLOCK_50) 
		begin	
			if rising_edge(CLOCK_50) then
				acc <= acc+1;
				if acc >= to_unsigned(499, 9) then
					acc <= to_unsigned(0,9);
				end if;
			end if;
			 case acc is
					when "000000000" => sinVal <= "10000000000000";
					when "000000001" => sinVal <= "10000001100110";
					when "000000010" => sinVal <= "10000011001101";
					when "000000011" => sinVal <= "10000100110100";
					when "000000100" => sinVal <= "10000110011011";
					when "000000101" => sinVal <= "10001000000010";
					when "000000110" => sinVal <= "10001001101001";
					when "000000111" => sinVal <= "10001011001111";
					when "000001000" => sinVal <= "10001100110110";
					when "000001001" => sinVal <= "10001110011100";
					when "000001010" => sinVal <= "10010000000010";
					when "000001011" => sinVal <= "10010001101000";
					when "000001100" => sinVal <= "10010011001110";
					when "000001101" => sinVal <= "10010100110100";
					when "000001110" => sinVal <= "10010110011001";
					when "000001111" => sinVal <= "10010111111110";
					when "000010000" => sinVal <= "10011001100011";
					when "000010001" => sinVal <= "10011011001000";
					when "000010010" => sinVal <= "10011100101101";
					when "000010011" => sinVal <= "10011110010001";
					when "000010100" => sinVal <= "10011111110101";
					when "000010101" => sinVal <= "10100001011000";
					when "000010110" => sinVal <= "10100010111011";
					when "000010111" => sinVal <= "10100100011110";
					when "000011000" => sinVal <= "10100110000001";
					when "000011001" => sinVal <= "10100111100011";
					when "000011010" => sinVal <= "10101001000101";
					when "000011011" => sinVal <= "10101010100110";
					when "000011100" => sinVal <= "10101100000111";
					when "000011101" => sinVal <= "10101101100111";
					when "000011110" => sinVal <= "10101111000111";
					when "000011111" => sinVal <= "10110000100110";
					when "000100000" => sinVal <= "10110010000101";
					when "000100001" => sinVal <= "10110011100100";
					when "000100010" => sinVal <= "10110101000010";
					when "000100011" => sinVal <= "10110110011111";
					when "000100100" => sinVal <= "10110111111100";
					when "000100101" => sinVal <= "10111001011000";
					when "000100110" => sinVal <= "10111010110100";
					when "000100111" => sinVal <= "10111100001111";
					when "000101000" => sinVal <= "10111101101010";
					when "000101001" => sinVal <= "10111111000100";
					when "000101010" => sinVal <= "11000000011101";
					when "000101011" => sinVal <= "11000001110110";
					when "000101100" => sinVal <= "11000011001101";
					when "000101101" => sinVal <= "11000100100101";
					when "000101110" => sinVal <= "11000101111011";
					when "000101111" => sinVal <= "11000111010001";
					when "000110000" => sinVal <= "11001000100110";
					when "000110001" => sinVal <= "11001001111011";
					when "000110010" => sinVal <= "11001011001110";
					when "000110011" => sinVal <= "11001100100001";
					when "000110100" => sinVal <= "11001101110011";
					when "000110101" => sinVal <= "11001111000101";
					when "000110110" => sinVal <= "11010000010101";
					when "000110111" => sinVal <= "11010001100101";
					when "000111000" => sinVal <= "11010010110100";
					when "000111001" => sinVal <= "11010100000010";
					when "000111010" => sinVal <= "11010101001111";
					when "000111011" => sinVal <= "11010110011011";
					when "000111100" => sinVal <= "11010111100111";
					when "000111101" => sinVal <= "11011000110010";
					when "000111110" => sinVal <= "11011001111011";
					when "000111111" => sinVal <= "11011011000100";
					when "001000000" => sinVal <= "11011100001100";
					when "001000001" => sinVal <= "11011101010011";
					when "001000010" => sinVal <= "11011110011001";
					when "001000011" => sinVal <= "11011111011110";
					when "001000100" => sinVal <= "11100000100010";
					when "001000101" => sinVal <= "11100001100101";
					when "001000110" => sinVal <= "11100010100111";
					when "001000111" => sinVal <= "11100011101000";
					when "001001000" => sinVal <= "11100100101000";
					when "001001001" => sinVal <= "11100101100111";
					when "001001010" => sinVal <= "11100110100110";
					when "001001011" => sinVal <= "11100111100011";
					when "001001100" => sinVal <= "11101000011111";
					when "001001101" => sinVal <= "11101001011001";
					when "001001110" => sinVal <= "11101010010011";
					when "001001111" => sinVal <= "11101011001100";
					when "001010000" => sinVal <= "11101100000100";
					when "001010001" => sinVal <= "11101100111010";
					when "001010010" => sinVal <= "11101101110000";
					when "001010011" => sinVal <= "11101110100100";
					when "001010100" => sinVal <= "11101111011000";
					when "001010101" => sinVal <= "11110000001010";
					when "001010110" => sinVal <= "11110000111011";
					when "001010111" => sinVal <= "11110001101011";
					when "001011000" => sinVal <= "11110010011001";
					when "001011001" => sinVal <= "11110011000111";
					when "001011010" => sinVal <= "11110011110011";
					when "001011011" => sinVal <= "11110100011111";
					when "001011100" => sinVal <= "11110101001001";
					when "001011101" => sinVal <= "11110101110010";
					when "001011110" => sinVal <= "11110110011001";
					when "001011111" => sinVal <= "11110111000000";
					when "001100000" => sinVal <= "11110111100101";
					when "001100001" => sinVal <= "11111000001001";
					when "001100010" => sinVal <= "11111000101100";
					when "001100011" => sinVal <= "11111001001110";
					when "001100100" => sinVal <= "11111001101110";
					when "001100101" => sinVal <= "11111010001101";
					when "001100110" => sinVal <= "11111010101011";
					when "001100111" => sinVal <= "11111011001000";
					when "001101000" => sinVal <= "11111011100011";
					when "001101001" => sinVal <= "11111011111110";
					when "001101010" => sinVal <= "11111100010111";
					when "001101011" => sinVal <= "11111100101110";
					when "001101100" => sinVal <= "11111101000101";
					when "001101101" => sinVal <= "11111101011010";
					when "001101110" => sinVal <= "11111101101110";
					when "001101111" => sinVal <= "11111110000001";
					when "001110000" => sinVal <= "11111110010010";
					when "001110001" => sinVal <= "11111110100010";
					when "001110010" => sinVal <= "11111110110001";
					when "001110011" => sinVal <= "11111110111110";
					when "001110100" => sinVal <= "11111111001011";
					when "001110101" => sinVal <= "11111111010110";
					when "001110110" => sinVal <= "11111111011111";
					when "001110111" => sinVal <= "11111111101000";
					when "001111000" => sinVal <= "11111111101111";
					when "001111001" => sinVal <= "11111111110101";
					when "001111010" => sinVal <= "11111111111001";
					when "001111011" => sinVal <= "11111111111100";
					when "001111100" => sinVal <= "11111111111110";
					when "001111101" => sinVal <= "11111111111111";
					when "001111110" => sinVal <= "11111111111110";
					when "001111111" => sinVal <= "11111111111100";
					when "010000000" => sinVal <= "11111111111001";
					when "010000001" => sinVal <= "11111111110101";
					when "010000010" => sinVal <= "11111111101111";
					when "010000011" => sinVal <= "11111111101000";
					when "010000100" => sinVal <= "11111111011111";
					when "010000101" => sinVal <= "11111111010110";
					when "010000110" => sinVal <= "11111111001011";
					when "010000111" => sinVal <= "11111110111110";
					when "010001000" => sinVal <= "11111110110001";
					when "010001001" => sinVal <= "11111110100010";
					when "010001010" => sinVal <= "11111110010010";
					when "010001011" => sinVal <= "11111110000001";
					when "010001100" => sinVal <= "11111101101110";
					when "010001101" => sinVal <= "11111101011010";
					when "010001110" => sinVal <= "11111101000101";
					when "010001111" => sinVal <= "11111100101110";
					when "010010000" => sinVal <= "11111100010111";
					when "010010001" => sinVal <= "11111011111110";
					when "010010010" => sinVal <= "11111011100011";
					when "010010011" => sinVal <= "11111011001000";
					when "010010100" => sinVal <= "11111010101011";
					when "010010101" => sinVal <= "11111010001101";
					when "010010110" => sinVal <= "11111001101110";
					when "010010111" => sinVal <= "11111001001110";
					when "010011000" => sinVal <= "11111000101100";
					when "010011001" => sinVal <= "11111000001001";
					when "010011010" => sinVal <= "11110111100101";
					when "010011011" => sinVal <= "11110111000000";
					when "010011100" => sinVal <= "11110110011001";
					when "010011101" => sinVal <= "11110101110010";
					when "010011110" => sinVal <= "11110101001001";
					when "010011111" => sinVal <= "11110100011111";
					when "010100000" => sinVal <= "11110011110011";
					when "010100001" => sinVal <= "11110011000111";
					when "010100010" => sinVal <= "11110010011001";
					when "010100011" => sinVal <= "11110001101011";
					when "010100100" => sinVal <= "11110000111011";
					when "010100101" => sinVal <= "11110000001010";
					when "010100110" => sinVal <= "11101111011000";
					when "010100111" => sinVal <= "11101110100100";
					when "010101000" => sinVal <= "11101101110000";
					when "010101001" => sinVal <= "11101100111010";
					when "010101010" => sinVal <= "11101100000100";
					when "010101011" => sinVal <= "11101011001100";
					when "010101100" => sinVal <= "11101010010011";
					when "010101101" => sinVal <= "11101001011001";
					when "010101110" => sinVal <= "11101000011111";
					when "010101111" => sinVal <= "11100111100011";
					when "010110000" => sinVal <= "11100110100110";
					when "010110001" => sinVal <= "11100101100111";
					when "010110010" => sinVal <= "11100100101000";
					when "010110011" => sinVal <= "11100011101000";
					when "010110100" => sinVal <= "11100010100111";
					when "010110101" => sinVal <= "11100001100101";
					when "010110110" => sinVal <= "11100000100010";
					when "010110111" => sinVal <= "11011111011110";
					when "010111000" => sinVal <= "11011110011001";
					when "010111001" => sinVal <= "11011101010011";
					when "010111010" => sinVal <= "11011100001100";
					when "010111011" => sinVal <= "11011011000100";
					when "010111100" => sinVal <= "11011001111011";
					when "010111101" => sinVal <= "11011000110010";
					when "010111110" => sinVal <= "11010111100111";
					when "010111111" => sinVal <= "11010110011011";
					when "011000000" => sinVal <= "11010101001111";
					when "011000001" => sinVal <= "11010100000010";
					when "011000010" => sinVal <= "11010010110100";
					when "011000011" => sinVal <= "11010001100101";
					when "011000100" => sinVal <= "11010000010101";
					when "011000101" => sinVal <= "11001111000101";
					when "011000110" => sinVal <= "11001101110011";
					when "011000111" => sinVal <= "11001100100001";
					when "011001000" => sinVal <= "11001011001110";
					when "011001001" => sinVal <= "11001001111011";
					when "011001010" => sinVal <= "11001000100110";
					when "011001011" => sinVal <= "11000111010001";
					when "011001100" => sinVal <= "11000101111011";
					when "011001101" => sinVal <= "11000100100101";
					when "011001110" => sinVal <= "11000011001101";
					when "011001111" => sinVal <= "11000001110110";
					when "011010000" => sinVal <= "11000000011101";
					when "011010001" => sinVal <= "10111111000100";
					when "011010010" => sinVal <= "10111101101010";
					when "011010011" => sinVal <= "10111100001111";
					when "011010100" => sinVal <= "10111010110100";
					when "011010101" => sinVal <= "10111001011000";
					when "011010110" => sinVal <= "10110111111100";
					when "011010111" => sinVal <= "10110110011111";
					when "011011000" => sinVal <= "10110101000010";
					when "011011001" => sinVal <= "10110011100100";
					when "011011010" => sinVal <= "10110010000101";
					when "011011011" => sinVal <= "10110000100110";
					when "011011100" => sinVal <= "10101111000111";
					when "011011101" => sinVal <= "10101101100111";
					when "011011110" => sinVal <= "10101100000111";
					when "011011111" => sinVal <= "10101010100110";
					when "011100000" => sinVal <= "10101001000101";
					when "011100001" => sinVal <= "10100111100011";
					when "011100010" => sinVal <= "10100110000001";
					when "011100011" => sinVal <= "10100100011110";
					when "011100100" => sinVal <= "10100010111011";
					when "011100101" => sinVal <= "10100001011000";
					when "011100110" => sinVal <= "10011111110101";
					when "011100111" => sinVal <= "10011110010001";
					when "011101000" => sinVal <= "10011100101101";
					when "011101001" => sinVal <= "10011011001000";
					when "011101010" => sinVal <= "10011001100011";
					when "011101011" => sinVal <= "10010111111110";
					when "011101100" => sinVal <= "10010110011001";
					when "011101101" => sinVal <= "10010100110100";
					when "011101110" => sinVal <= "10010011001110";
					when "011101111" => sinVal <= "10010001101000";
					when "011110000" => sinVal <= "10010000000010";
					when "011110001" => sinVal <= "10001110011100";
					when "011110010" => sinVal <= "10001100110110";
					when "011110011" => sinVal <= "10001011001111";
					when "011110100" => sinVal <= "10001001101001";
					when "011110101" => sinVal <= "10001000000010";
					when "011110110" => sinVal <= "10000110011011";
					when "011110111" => sinVal <= "10000100110100";
					when "011111000" => sinVal <= "10000011001101";
					when "011111001" => sinVal <= "10000001100110";
					when "011111010" => sinVal <= "10000000000000";
					when "011111011" => sinVal <= "01111110011001";
					when "011111100" => sinVal <= "01111100110010";
					when "011111101" => sinVal <= "01111011001011";
					when "011111110" => sinVal <= "01111001100100";
					when "011111111" => sinVal <= "01110111111101";
					when "100000000" => sinVal <= "01110110010110";
					when "100000001" => sinVal <= "01110100110000";
					when "100000010" => sinVal <= "01110011001001";
					when "100000011" => sinVal <= "01110001100011";
					when "100000100" => sinVal <= "01101111111101";
					when "100000101" => sinVal <= "01101110010111";
					when "100000110" => sinVal <= "01101100110001";
					when "100000111" => sinVal <= "01101011001011";
					when "100001000" => sinVal <= "01101001100110";
					when "100001001" => sinVal <= "01101000000001";
					when "100001010" => sinVal <= "01100110011100";
					when "100001011" => sinVal <= "01100100110111";
					when "100001100" => sinVal <= "01100011010010";
					when "100001101" => sinVal <= "01100001101110";
					when "100001110" => sinVal <= "01100000001010";
					when "100001111" => sinVal <= "01011110100111";
					when "100010000" => sinVal <= "01011101000100";
					when "100010001" => sinVal <= "01011011100001";
					when "100010010" => sinVal <= "01011001111110";
					when "100010011" => sinVal <= "01011000011100";
					when "100010100" => sinVal <= "01010110111010";
					when "100010101" => sinVal <= "01010101011001";
					when "100010110" => sinVal <= "01010011111000";
					when "100010111" => sinVal <= "01010010011000";
					when "100011000" => sinVal <= "01010000111000";
					when "100011001" => sinVal <= "01001111011001";
					when "100011010" => sinVal <= "01001101111010";
					when "100011011" => sinVal <= "01001100011011";
					when "100011100" => sinVal <= "01001010111101";
					when "100011101" => sinVal <= "01001001100000";
					when "100011110" => sinVal <= "01001000000011";
					when "100011111" => sinVal <= "01000110100111";
					when "100100000" => sinVal <= "01000101001011";
					when "100100001" => sinVal <= "01000011110000";
					when "100100010" => sinVal <= "01000010010101";
					when "100100011" => sinVal <= "01000000111011";
					when "100100100" => sinVal <= "00111111100010";
					when "100100101" => sinVal <= "00111110001001";
					when "100100110" => sinVal <= "00111100110010";
					when "100100111" => sinVal <= "00111011011010";
					when "100101000" => sinVal <= "00111010000100";
					when "100101001" => sinVal <= "00111000101110";
					when "100101010" => sinVal <= "00110111011001";
					when "100101011" => sinVal <= "00110110000100";
					when "100101100" => sinVal <= "00110100110001";
					when "100101101" => sinVal <= "00110011011110";
					when "100101110" => sinVal <= "00110010001100";
					when "100101111" => sinVal <= "00110000111010";
					when "100110000" => sinVal <= "00101111101010";
					when "100110001" => sinVal <= "00101110011010";
					when "100110010" => sinVal <= "00101101001011";
					when "100110011" => sinVal <= "00101011111101";
					when "100110100" => sinVal <= "00101010110000";
					when "100110101" => sinVal <= "00101001100100";
					when "100110110" => sinVal <= "00101000011000";
					when "100110111" => sinVal <= "00100111001101";
					when "100111000" => sinVal <= "00100110000100";
					when "100111001" => sinVal <= "00100100111011";
					when "100111010" => sinVal <= "00100011110011";
					when "100111011" => sinVal <= "00100010101100";
					when "100111100" => sinVal <= "00100001100110";
					when "100111101" => sinVal <= "00100000100001";
					when "100111110" => sinVal <= "00011111011101";
					when "100111111" => sinVal <= "00011110011010";
					when "101000000" => sinVal <= "00011101011000";
					when "101000001" => sinVal <= "00011100010111";
					when "101000010" => sinVal <= "00011011010111";
					when "101000011" => sinVal <= "00011010011000";
					when "101000100" => sinVal <= "00011001011001";
					when "101000101" => sinVal <= "00011000011100";
					when "101000110" => sinVal <= "00010111100000";
					when "101000111" => sinVal <= "00010110100110";
					when "101001000" => sinVal <= "00010101101100";
					when "101001001" => sinVal <= "00010100110011";
					when "101001010" => sinVal <= "00010011111011";
					when "101001011" => sinVal <= "00010011000101";
					when "101001100" => sinVal <= "00010010001111";
					when "101001101" => sinVal <= "00010001011011";
					when "101001110" => sinVal <= "00010000100111";
					when "101001111" => sinVal <= "00001111110101";
					when "101010000" => sinVal <= "00001111000100";
					when "101010001" => sinVal <= "00001110010100";
					when "101010010" => sinVal <= "00001101100110";
					when "101010011" => sinVal <= "00001100111000";
					when "101010100" => sinVal <= "00001100001100";
					when "101010101" => sinVal <= "00001011100000";
					when "101010110" => sinVal <= "00001010110110";
					when "101010111" => sinVal <= "00001010001101";
					when "101011000" => sinVal <= "00001001100110";
					when "101011001" => sinVal <= "00001000111111";
					when "101011010" => sinVal <= "00001000011010";
					when "101011011" => sinVal <= "00000111110110";
					when "101011100" => sinVal <= "00000111010011";
					when "101011101" => sinVal <= "00000110110001";
					when "101011110" => sinVal <= "00000110010001";
					when "101011111" => sinVal <= "00000101110010";
					when "101100000" => sinVal <= "00000101010100";
					when "101100001" => sinVal <= "00000100110111";
					when "101100010" => sinVal <= "00000100011100";
					when "101100011" => sinVal <= "00000100000001";
					when "101100100" => sinVal <= "00000011101000";
					when "101100101" => sinVal <= "00000011010001";
					when "101100110" => sinVal <= "00000010111010";
					when "101100111" => sinVal <= "00000010100101";
					when "101101000" => sinVal <= "00000010010001";
					when "101101001" => sinVal <= "00000001111110";
					when "101101010" => sinVal <= "00000001101101";
					when "101101011" => sinVal <= "00000001011101";
					when "101101100" => sinVal <= "00000001001110";
					when "101101101" => sinVal <= "00000001000001";
					when "101101110" => sinVal <= "00000000110100";
					when "101101111" => sinVal <= "00000000101001";
					when "101110000" => sinVal <= "00000000100000";
					when "101110001" => sinVal <= "00000000010111";
					when "101110010" => sinVal <= "00000000010000";
					when "101110011" => sinVal <= "00000000001010";
					when "101110100" => sinVal <= "00000000000110";
					when "101110101" => sinVal <= "00000000000011";
					when "101110110" => sinVal <= "00000000000001";
					when "101110111" => sinVal <= "00000000000000";
					when "101111000" => sinVal <= "00000000000001";
					when "101111001" => sinVal <= "00000000000011";
					when "101111010" => sinVal <= "00000000000110";
					when "101111011" => sinVal <= "00000000001010";
					when "101111100" => sinVal <= "00000000010000";
					when "101111101" => sinVal <= "00000000010111";
					when "101111110" => sinVal <= "00000000100000";
					when "101111111" => sinVal <= "00000000101001";
					when "110000000" => sinVal <= "00000000110100";
					when "110000001" => sinVal <= "00000001000001";
					when "110000010" => sinVal <= "00000001001110";
					when "110000011" => sinVal <= "00000001011101";
					when "110000100" => sinVal <= "00000001101101";
					when "110000101" => sinVal <= "00000001111110";
					when "110000110" => sinVal <= "00000010010001";
					when "110000111" => sinVal <= "00000010100101";
					when "110001000" => sinVal <= "00000010111010";
					when "110001001" => sinVal <= "00000011010001";
					when "110001010" => sinVal <= "00000011101000";
					when "110001011" => sinVal <= "00000100000001";
					when "110001100" => sinVal <= "00000100011100";
					when "110001101" => sinVal <= "00000100110111";
					when "110001110" => sinVal <= "00000101010100";
					when "110001111" => sinVal <= "00000101110010";
					when "110010000" => sinVal <= "00000110010001";
					when "110010001" => sinVal <= "00000110110001";
					when "110010010" => sinVal <= "00000111010011";
					when "110010011" => sinVal <= "00000111110110";
					when "110010100" => sinVal <= "00001000011010";
					when "110010101" => sinVal <= "00001000111111";
					when "110010110" => sinVal <= "00001001100110";
					when "110010111" => sinVal <= "00001010001101";
					when "110011000" => sinVal <= "00001010110110";
					when "110011001" => sinVal <= "00001011100000";
					when "110011010" => sinVal <= "00001100001100";
					when "110011011" => sinVal <= "00001100111000";
					when "110011100" => sinVal <= "00001101100110";
					when "110011101" => sinVal <= "00001110010100";
					when "110011110" => sinVal <= "00001111000100";
					when "110011111" => sinVal <= "00001111110101";
					when "110100000" => sinVal <= "00010000100111";
					when "110100001" => sinVal <= "00010001011011";
					when "110100010" => sinVal <= "00010010001111";
					when "110100011" => sinVal <= "00010011000101";
					when "110100100" => sinVal <= "00010011111011";
					when "110100101" => sinVal <= "00010100110011";
					when "110100110" => sinVal <= "00010101101100";
					when "110100111" => sinVal <= "00010110100110";
					when "110101000" => sinVal <= "00010111100000";
					when "110101001" => sinVal <= "00011000011100";
					when "110101010" => sinVal <= "00011001011001";
					when "110101011" => sinVal <= "00011010011000";
					when "110101100" => sinVal <= "00011011010111";
					when "110101101" => sinVal <= "00011100010111";
					when "110101110" => sinVal <= "00011101011000";
					when "110101111" => sinVal <= "00011110011010";
					when "110110000" => sinVal <= "00011111011101";
					when "110110001" => sinVal <= "00100000100001";
					when "110110010" => sinVal <= "00100001100110";
					when "110110011" => sinVal <= "00100010101100";
					when "110110100" => sinVal <= "00100011110011";
					when "110110101" => sinVal <= "00100100111011";
					when "110110110" => sinVal <= "00100110000100";
					when "110110111" => sinVal <= "00100111001101";
					when "110111000" => sinVal <= "00101000011000";
					when "110111001" => sinVal <= "00101001100100";
					when "110111010" => sinVal <= "00101010110000";
					when "110111011" => sinVal <= "00101011111101";
					when "110111100" => sinVal <= "00101101001011";
					when "110111101" => sinVal <= "00101110011010";
					when "110111110" => sinVal <= "00101111101010";
					when "110111111" => sinVal <= "00110000111010";
					when "111000000" => sinVal <= "00110010001100";
					when "111000001" => sinVal <= "00110011011110";
					when "111000010" => sinVal <= "00110100110001";
					when "111000011" => sinVal <= "00110110000100";
					when "111000100" => sinVal <= "00110111011001";
					when "111000101" => sinVal <= "00111000101110";
					when "111000110" => sinVal <= "00111010000100";
					when "111000111" => sinVal <= "00111011011010";
					when "111001000" => sinVal <= "00111100110010";
					when "111001001" => sinVal <= "00111110001001";
					when "111001010" => sinVal <= "00111111100010";
					when "111001011" => sinVal <= "01000000111011";
					when "111001100" => sinVal <= "01000010010101";
					when "111001101" => sinVal <= "01000011110000";
					when "111001110" => sinVal <= "01000101001011";
					when "111001111" => sinVal <= "01000110100111";
					when "111010000" => sinVal <= "01001000000011";
					when "111010001" => sinVal <= "01001001100000";
					when "111010010" => sinVal <= "01001010111101";
					when "111010011" => sinVal <= "01001100011011";
					when "111010100" => sinVal <= "01001101111010";
					when "111010101" => sinVal <= "01001111011001";
					when "111010110" => sinVal <= "01010000111000";
					when "111010111" => sinVal <= "01010010011000";
					when "111011000" => sinVal <= "01010011111000";
					when "111011001" => sinVal <= "01010101011001";
					when "111011010" => sinVal <= "01010110111010";
					when "111011011" => sinVal <= "01011000011100";
					when "111011100" => sinVal <= "01011001111110";
					when "111011101" => sinVal <= "01011011100001";
					when "111011110" => sinVal <= "01011101000100";
					when "111011111" => sinVal <= "01011110100111";
					when "111100000" => sinVal <= "01100000001010";
					when "111100001" => sinVal <= "01100001101110";
					when "111100010" => sinVal <= "01100011010010";
					when "111100011" => sinVal <= "01100100110111";
					when "111100100" => sinVal <= "01100110011100";
					when "111100101" => sinVal <= "01101000000001";
					when "111100110" => sinVal <= "01101001100110";
					when "111100111" => sinVal <= "01101011001011";
					when "111101000" => sinVal <= "01101100110001";
					when "111101001" => sinVal <= "01101110010111";
					when "111101010" => sinVal <= "01101111111101";
					when "111101011" => sinVal <= "01110001100011";
					when "111101100" => sinVal <= "01110011001001";
					when "111101101" => sinVal <= "01110100110000";
					when "111101110" => sinVal <= "01110110010110";
					when "111101111" => sinVal <= "01110111111101";
					when "111110000" => sinVal <= "01111001100100";
					when "111110001" => sinVal <= "01111011001011";
					when "111110010" => sinVal <= "01111100110010";
					when "111110011" => sinVal <= "01111110011001";
					when others => sinVal <= "00000000000000";
				 end case;
	end process; 
	
	audio1: DE2_Audio_Example port map(sinVal, CLOCK_50, CLOCK_27, KEY, AUD_ADCDAT, 
	AUD_BCLK, AUD_ADCLRCK, AUD_DACLRCK, I2C_SDAT, AUD_XCK, AUD_DACDAT, I2C_SCLK, LEDR, SW);
end architecture behaviour;