
module nios_system2 (
	audio_ADCDAT,
	audio_ADCLRCK,
	audio_BCLK,
	audio_DACDAT,
	audio_DACLRCK,
	audio_clk_clk,
	audio_irq_irq,
	audio_pll_ref_clk_clk,
	audio_pll_ref_reset_reset,
	audio_reset_reset,
	audio_slave_address,
	audio_slave_chipselect,
	audio_slave_read,
	audio_slave_write,
	audio_slave_writedata,
	audio_slave_readdata,
	av_config_SDAT,
	av_config_SCLK,
	clk_clk,
	expansion_jp5_export,
	flash_ADDR,
	flash_CE_N,
	flash_OE_N,
	flash_WE_N,
	flash_RST_N,
	flash_DQ,
	green_leds_export,
	pushbuttons_export,
	red_leds_export,
	reset_reset_n,
	sdram_addr,
	sdram_ba,
	sdram_cas_n,
	sdram_cke,
	sdram_cs_n,
	sdram_dq,
	sdram_dqm,
	sdram_ras_n,
	sdram_we_n,
	serial_port_RXD,
	serial_port_TXD,
	slider_switches_export,
	sram_DQ,
	sram_ADDR,
	sram_LB_N,
	sram_UB_N,
	sram_CE_N,
	sram_OE_N,
	sram_WE_N,
	video_ext_PIXEL_CLK,
	video_ext_LINE_VALID,
	video_ext_FRAME_VALID,
	video_ext_pixel_clk_reset,
	video_ext_PIXEL_DATA);	

	input		audio_ADCDAT;
	input		audio_ADCLRCK;
	input		audio_BCLK;
	output		audio_DACDAT;
	input		audio_DACLRCK;
	output		audio_clk_clk;
	output		audio_irq_irq;
	input		audio_pll_ref_clk_clk;
	input		audio_pll_ref_reset_reset;
	output		audio_reset_reset;
	input	[1:0]	audio_slave_address;
	input		audio_slave_chipselect;
	input		audio_slave_read;
	input		audio_slave_write;
	input	[31:0]	audio_slave_writedata;
	output	[31:0]	audio_slave_readdata;
	inout		av_config_SDAT;
	output		av_config_SCLK;
	input		clk_clk;
	inout	[31:0]	expansion_jp5_export;
	output	[22:0]	flash_ADDR;
	output		flash_CE_N;
	output		flash_OE_N;
	output		flash_WE_N;
	output		flash_RST_N;
	inout	[7:0]	flash_DQ;
	output	[8:0]	green_leds_export;
	input	[3:0]	pushbuttons_export;
	output	[17:0]	red_leds_export;
	input		reset_reset_n;
	output	[12:0]	sdram_addr;
	output	[1:0]	sdram_ba;
	output		sdram_cas_n;
	output		sdram_cke;
	output		sdram_cs_n;
	inout	[31:0]	sdram_dq;
	output	[3:0]	sdram_dqm;
	output		sdram_ras_n;
	output		sdram_we_n;
	input		serial_port_RXD;
	output		serial_port_TXD;
	input	[17:0]	slider_switches_export;
	inout	[15:0]	sram_DQ;
	output	[19:0]	sram_ADDR;
	output		sram_LB_N;
	output		sram_UB_N;
	output		sram_CE_N;
	output		sram_OE_N;
	output		sram_WE_N;
	input		video_ext_PIXEL_CLK;
	input		video_ext_LINE_VALID;
	input		video_ext_FRAME_VALID;
	input		video_ext_pixel_clk_reset;
	input	[11:0]	video_ext_PIXEL_DATA;
endmodule
