-- nios_system.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_system is
	port (
		audio_ADCDAT                : in    std_logic                     := '0';             --                audio.ADCDAT
		audio_ADCLRCK               : in    std_logic                     := '0';             --                     .ADCLRCK
		audio_BCLK                  : in    std_logic                     := '0';             --                     .BCLK
		audio_DACDAT                : out   std_logic;                                        --                     .DACDAT
		audio_DACLRCK               : in    std_logic                     := '0';             --                     .DACLRCK
		audio_clk_clk               : out   std_logic;                                        --            audio_clk.clk
		audio_pll_ref_clk_clk       : in    std_logic                     := '0';             --    audio_pll_ref_clk.clk
		audio_pll_ref_reset_reset   : in    std_logic                     := '0';             --  audio_pll_ref_reset.reset
		av_config_SDAT              : inout std_logic                     := '0';             --            av_config.SDAT
		av_config_SCLK              : out   std_logic;                                        --                     .SCLK
		expansion_jp5_export        : inout std_logic_vector(31 downto 0) := (others => '0'); --        expansion_jp5.export
		flash_ADDR                  : out   std_logic_vector(22 downto 0);                    --                flash.ADDR
		flash_CE_N                  : out   std_logic;                                        --                     .CE_N
		flash_OE_N                  : out   std_logic;                                        --                     .OE_N
		flash_WE_N                  : out   std_logic;                                        --                     .WE_N
		flash_RST_N                 : out   std_logic;                                        --                     .RST_N
		flash_DQ                    : inout std_logic_vector(7 downto 0)  := (others => '0'); --                     .DQ
		green_leds_export           : out   std_logic_vector(8 downto 0);                     --           green_leds.export
		pushbuttons_export          : in    std_logic_vector(3 downto 0)  := (others => '0'); --          pushbuttons.export
		red_leds_export             : out   std_logic_vector(17 downto 0);                    --             red_leds.export
		sdram_addr                  : out   std_logic_vector(12 downto 0);                    --                sdram.addr
		sdram_ba                    : out   std_logic_vector(1 downto 0);                     --                     .ba
		sdram_cas_n                 : out   std_logic;                                        --                     .cas_n
		sdram_cke                   : out   std_logic;                                        --                     .cke
		sdram_cs_n                  : out   std_logic;                                        --                     .cs_n
		sdram_dq                    : inout std_logic_vector(31 downto 0) := (others => '0'); --                     .dq
		sdram_dqm                   : out   std_logic_vector(3 downto 0);                     --                     .dqm
		sdram_ras_n                 : out   std_logic;                                        --                     .ras_n
		sdram_we_n                  : out   std_logic;                                        --                     .we_n
		sdram_clk_clk               : out   std_logic;                                        --            sdram_clk.clk
		serial_port_RXD             : in    std_logic                     := '0';             --          serial_port.RXD
		serial_port_TXD             : out   std_logic;                                        --                     .TXD
		slider_switches_export      : in    std_logic_vector(17 downto 0) := (others => '0'); --      slider_switches.export
		sram_DQ                     : inout std_logic_vector(15 downto 0) := (others => '0'); --                 sram.DQ
		sram_ADDR                   : out   std_logic_vector(19 downto 0);                    --                     .ADDR
		sram_LB_N                   : out   std_logic;                                        --                     .LB_N
		sram_UB_N                   : out   std_logic;                                        --                     .UB_N
		sram_CE_N                   : out   std_logic;                                        --                     .CE_N
		sram_OE_N                   : out   std_logic;                                        --                     .OE_N
		sram_WE_N                   : out   std_logic;                                        --                     .WE_N
		system_pll_ref_clk_clk      : in    std_logic                     := '0';             --   system_pll_ref_clk.clk
		system_pll_ref_reset_reset  : in    std_logic                     := '0';             -- system_pll_ref_reset.reset
		video_ext_1_PIXEL_CLK       : in    std_logic                     := '0';             --          video_ext_1.PIXEL_CLK
		video_ext_1_LINE_VALID      : in    std_logic                     := '0';             --                     .LINE_VALID
		video_ext_1_FRAME_VALID     : in    std_logic                     := '0';             --                     .FRAME_VALID
		video_ext_1_pixel_clk_reset : in    std_logic                     := '0';             --                     .pixel_clk_reset
		video_ext_1_PIXEL_DATA      : in    std_logic_vector(11 downto 0) := (others => '0')  --                     .PIXEL_DATA
	);
end entity nios_system;

architecture rtl of nios_system is
	component nios_system_AV_Config is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component nios_system_AV_Config;

	component nios_system_Audio_Subsystem is
		port (
			audio_ADCDAT              : in  std_logic                     := 'X';             -- ADCDAT
			audio_ADCLRCK             : in  std_logic                     := 'X';             -- ADCLRCK
			audio_BCLK                : in  std_logic                     := 'X';             -- BCLK
			audio_DACDAT              : out std_logic;                                        -- DACDAT
			audio_DACLRCK             : in  std_logic                     := 'X';             -- DACLRCK
			audio_clk_clk             : out std_logic;                                        -- clk
			audio_irq_irq             : out std_logic;                                        -- irq
			audio_pll_ref_clk_clk     : in  std_logic                     := 'X';             -- clk
			audio_pll_ref_reset_reset : in  std_logic                     := 'X';             -- reset
			audio_reset_reset         : out std_logic;                                        -- reset
			audio_slave_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			audio_slave_chipselect    : in  std_logic                     := 'X';             -- chipselect
			audio_slave_read          : in  std_logic                     := 'X';             -- read
			audio_slave_write         : in  std_logic                     := 'X';             -- write
			audio_slave_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			audio_slave_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			sys_clk_clk               : in  std_logic                     := 'X';             -- clk
			sys_reset_reset_n         : in  std_logic                     := 'X'              -- reset_n
		);
	end component nios_system_Audio_Subsystem;

	component nios_system_CameraD5M_0 is
		port (
			camera_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			clk_clk                   : in  std_logic                     := 'X';             -- clk
			reset_reset_n             : in  std_logic                     := 'X';             -- reset_n
			video_ext_PIXEL_CLK       : in  std_logic                     := 'X';             -- PIXEL_CLK
			video_ext_LINE_VALID      : in  std_logic                     := 'X';             -- LINE_VALID
			video_ext_FRAME_VALID     : in  std_logic                     := 'X';             -- FRAME_VALID
			video_ext_pixel_clk_reset : in  std_logic                     := 'X';             -- pixel_clk_reset
			video_ext_PIXEL_DATA      : in  std_logic_vector(11 downto 0) := (others => 'X')  -- PIXEL_DATA
		);
	end component nios_system_CameraD5M_0;

	component nios_system_Expansion_JP5 is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset      : in    std_logic                     := 'X';             -- reset
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in    std_logic                     := 'X';             -- chipselect
			read       : in    std_logic                     := 'X';             -- read
			write      : in    std_logic                     := 'X';             -- write
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			GPIO       : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			irq        : out   std_logic                                         -- irq
		);
	end component nios_system_Expansion_JP5;

	component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface is
		generic (
			FLASH_MEMORY_ADDRESS_WIDTH : integer := 22
		);
		port (
			i_avalon_chip_select       : in    std_logic                     := 'X';             -- chipselect
			i_avalon_write             : in    std_logic                     := 'X';             -- write
			i_avalon_read              : in    std_logic                     := 'X';             -- read
			i_avalon_address           : in    std_logic_vector(20 downto 0) := (others => 'X'); -- address
			i_avalon_byteenable        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_avalon_writedata         : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			o_avalon_readdata          : out   std_logic_vector(31 downto 0);                    -- readdata
			o_avalon_waitrequest       : out   std_logic;                                        -- waitrequest
			i_clock                    : in    std_logic                     := 'X';             -- clk
			i_reset_n                  : in    std_logic                     := 'X';             -- reset_n
			FL_ADDR                    : out   std_logic_vector(22 downto 0);                    -- export
			FL_CE_N                    : out   std_logic;                                        -- export
			FL_OE_N                    : out   std_logic;                                        -- export
			FL_WE_N                    : out   std_logic;                                        -- export
			FL_RST_N                   : out   std_logic;                                        -- export
			FL_DQ                      : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			i_avalon_erase_write       : in    std_logic                     := 'X';             -- write
			i_avalon_erase_read        : in    std_logic                     := 'X';             -- read
			i_avalon_erase_byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_avalon_erase_writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			i_avalon_erase_chip_select : in    std_logic                     := 'X';             -- chipselect
			o_avalon_erase_readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			o_avalon_erase_waitrequest : out   std_logic                                         -- waitrequest
		);
	end component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface;

	component nios_system_Green_LEDs is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			LEDG       : out std_logic_vector(8 downto 0)                      -- export
		);
	end component nios_system_Green_LEDs;

	component nios_system_Interval_Timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_system_Interval_Timer;

	component nios_system_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_system_JTAG_UART;

	component nios_system_JTAG_to_FPGA_Bridge is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component nios_system_JTAG_to_FPGA_Bridge;

	component fpoint_wrapper is
		generic (
			useDivider : integer := 0
		);
		port (
			clk    : in  std_logic                     := 'X';             -- clk
			clk_en : in  std_logic                     := 'X';             -- clk_en
			dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			n      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- n
			reset  : in  std_logic                     := 'X';             -- reset
			start  : in  std_logic                     := 'X';             -- start
			done   : out std_logic;                                        -- done
			result : out std_logic_vector(31 downto 0)                     -- result
		);
	end component fpoint_wrapper;

	component nios_system_Processor1 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			E_ci_multi_done                     : in  std_logic                     := 'X';             -- done
			E_ci_multi_clk_en                   : out std_logic;                                        -- clk_en
			E_ci_multi_start                    : out std_logic;                                        -- start
			E_ci_result                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			D_ci_a                              : out std_logic_vector(4 downto 0);                     -- a
			D_ci_b                              : out std_logic_vector(4 downto 0);                     -- b
			D_ci_c                              : out std_logic_vector(4 downto 0);                     -- c
			D_ci_n                              : out std_logic_vector(7 downto 0);                     -- n
			D_ci_readra                         : out std_logic;                                        -- readra
			D_ci_readrb                         : out std_logic;                                        -- readrb
			D_ci_writerc                        : out std_logic;                                        -- writerc
			E_ci_dataa                          : out std_logic_vector(31 downto 0);                    -- dataa
			E_ci_datab                          : out std_logic_vector(31 downto 0);                    -- datab
			E_ci_multi_clock                    : out std_logic;                                        -- clk
			E_ci_multi_reset                    : out std_logic;                                        -- reset
			E_ci_multi_reset_req                : out std_logic;                                        -- reset_req
			W_ci_estatus                        : out std_logic;                                        -- estatus
			W_ci_ipending                       : out std_logic_vector(31 downto 0)                     -- ipending
		);
	end component nios_system_Processor1;

	component nios_system_Processor2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			E_ci_multi_done                     : in  std_logic                     := 'X';             -- done
			E_ci_multi_clk_en                   : out std_logic;                                        -- clk_en
			E_ci_multi_start                    : out std_logic;                                        -- start
			E_ci_result                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			D_ci_a                              : out std_logic_vector(4 downto 0);                     -- a
			D_ci_b                              : out std_logic_vector(4 downto 0);                     -- b
			D_ci_c                              : out std_logic_vector(4 downto 0);                     -- c
			D_ci_n                              : out std_logic_vector(7 downto 0);                     -- n
			D_ci_readra                         : out std_logic;                                        -- readra
			D_ci_readrb                         : out std_logic;                                        -- readrb
			D_ci_writerc                        : out std_logic;                                        -- writerc
			E_ci_dataa                          : out std_logic_vector(31 downto 0);                    -- dataa
			E_ci_datab                          : out std_logic_vector(31 downto 0);                    -- datab
			E_ci_multi_clock                    : out std_logic;                                        -- clk
			E_ci_multi_reset                    : out std_logic;                                        -- reset
			E_ci_multi_reset_req                : out std_logic;                                        -- reset_req
			W_ci_estatus                        : out std_logic;                                        -- estatus
			W_ci_ipending                       : out std_logic_vector(31 downto 0)                     -- ipending
		);
	end component nios_system_Processor2;

	component nios_system_Pushbuttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			KEY        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios_system_Pushbuttons;

	component nios_system_Red_LEDs is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			LEDR       : out std_logic_vector(17 downto 0)                     -- export
		);
	end component nios_system_Red_LEDs;

	component nios_system_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component nios_system_SDRAM;

	component nios_system_SRAM is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component nios_system_SRAM;

	component nios_system_Serial_Port is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic                     := 'X';             -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			irq        : out std_logic;                                        -- irq
			UART_RXD   : in  std_logic                     := 'X';             -- export
			UART_TXD   : out std_logic                                         -- export
		);
	end component nios_system_Serial_Port;

	component nios_system_Slider_Switches is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			SW         : in  std_logic_vector(17 downto 0) := (others => 'X')  -- export
		);
	end component nios_system_Slider_Switches;

	component nios_system_SysID is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios_system_SysID;

	component nios_system_System_PLL is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component nios_system_System_PLL;

	component altera_customins_master_translator is
		generic (
			SHARED_COMB_AND_MULTI : integer := 0
		);
		port (
			ci_slave_dataa            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result           : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra           : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb           : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc          : in  std_logic                     := 'X';             -- writerc
			ci_slave_a                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus          : in  std_logic                     := 'X';             -- estatus
			ci_slave_multi_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_multi_start      : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done       : out std_logic;                                        -- done
			comb_ci_master_dataa      : out std_logic_vector(31 downto 0);                    -- dataa
			comb_ci_master_datab      : out std_logic_vector(31 downto 0);                    -- datab
			comb_ci_master_result     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			comb_ci_master_n          : out std_logic_vector(7 downto 0);                     -- n
			comb_ci_master_readra     : out std_logic;                                        -- readra
			comb_ci_master_readrb     : out std_logic;                                        -- readrb
			comb_ci_master_writerc    : out std_logic;                                        -- writerc
			comb_ci_master_a          : out std_logic_vector(4 downto 0);                     -- a
			comb_ci_master_b          : out std_logic_vector(4 downto 0);                     -- b
			comb_ci_master_c          : out std_logic_vector(4 downto 0);                     -- c
			comb_ci_master_ipending   : out std_logic_vector(31 downto 0);                    -- ipending
			comb_ci_master_estatus    : out std_logic;                                        -- estatus
			multi_ci_master_clk       : out std_logic;                                        -- clk
			multi_ci_master_reset     : out std_logic;                                        -- reset
			multi_ci_master_clken     : out std_logic;                                        -- clk_en
			multi_ci_master_reset_req : out std_logic;                                        -- reset_req
			multi_ci_master_start     : out std_logic;                                        -- start
			multi_ci_master_done      : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra    : out std_logic;                                        -- readra
			multi_ci_master_readrb    : out std_logic;                                        -- readrb
			multi_ci_master_writerc   : out std_logic;                                        -- writerc
			multi_ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_slave_multi_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result     : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra     : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb     : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc    : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c          : in  std_logic_vector(4 downto 0)  := (others => 'X')  -- multi_c
		);
	end component altera_customins_master_translator;

	component nios_system_Processor1_custom_instruction_master_multi_xconnect is
		port (
			ci_slave_dataa       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result      : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra      : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb      : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc     : in  std_logic                     := 'X';             -- writerc
			ci_slave_a           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus     : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk         : in  std_logic                     := 'X';             -- clk
			ci_slave_reset       : in  std_logic                     := 'X';             -- reset
			ci_slave_clken       : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req   : in  std_logic                     := 'X';             -- reset_req
			ci_slave_start       : in  std_logic                     := 'X';             -- start
			ci_slave_done        : out std_logic;                                        -- done
			ci_master0_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n         : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra    : out std_logic;                                        -- readra
			ci_master0_readrb    : out std_logic;                                        -- readrb
			ci_master0_writerc   : out std_logic;                                        -- writerc
			ci_master0_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus   : out std_logic;                                        -- estatus
			ci_master0_clk       : out std_logic;                                        -- clk
			ci_master0_reset     : out std_logic;                                        -- reset
			ci_master0_clken     : out std_logic;                                        -- clk_en
			ci_master0_reset_req : out std_logic;                                        -- reset_req
			ci_master0_start     : out std_logic;                                        -- start
			ci_master0_done      : in  std_logic                     := 'X'              -- done
		);
	end component nios_system_Processor1_custom_instruction_master_multi_xconnect;

	component altera_customins_slave_translator is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_start      : in  std_logic                     := 'X';             -- start
			ci_slave_done       : out std_logic;                                        -- done
			ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master_n         : out std_logic_vector(1 downto 0);                     -- n
			ci_master_clk       : out std_logic;                                        -- clk
			ci_master_clken     : out std_logic;                                        -- clk_en
			ci_master_reset     : out std_logic;                                        -- reset
			ci_master_start     : out std_logic;                                        -- start
			ci_master_done      : in  std_logic                     := 'X';             -- done
			ci_master_readra    : out std_logic;                                        -- readra
			ci_master_readrb    : out std_logic;                                        -- readrb
			ci_master_writerc   : out std_logic;                                        -- writerc
			ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master_estatus   : out std_logic;                                        -- estatus
			ci_master_reset_req : out std_logic                                         -- reset_req
		);
	end component altera_customins_slave_translator;

	component nios_system_mm_interconnect_0 is
		port (
			System_PLL_sys_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			JTAG_UART_2nd_Core_reset_reset_bridge_in_reset_reset      : in  std_logic                     := 'X';             -- reset
			Processor1_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			Processor2_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			JTAG_to_FPGA_Bridge_master_address                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			JTAG_to_FPGA_Bridge_master_waitrequest                    : out std_logic;                                        -- waitrequest
			JTAG_to_FPGA_Bridge_master_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			JTAG_to_FPGA_Bridge_master_read                           : in  std_logic                     := 'X';             -- read
			JTAG_to_FPGA_Bridge_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			JTAG_to_FPGA_Bridge_master_readdatavalid                  : out std_logic;                                        -- readdatavalid
			JTAG_to_FPGA_Bridge_master_write                          : in  std_logic                     := 'X';             -- write
			JTAG_to_FPGA_Bridge_master_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Processor1_data_master_address                            : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			Processor1_data_master_waitrequest                        : out std_logic;                                        -- waitrequest
			Processor1_data_master_byteenable                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Processor1_data_master_read                               : in  std_logic                     := 'X';             -- read
			Processor1_data_master_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			Processor1_data_master_write                              : in  std_logic                     := 'X';             -- write
			Processor1_data_master_writedata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Processor1_data_master_debugaccess                        : in  std_logic                     := 'X';             -- debugaccess
			Processor1_instruction_master_address                     : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			Processor1_instruction_master_waitrequest                 : out std_logic;                                        -- waitrequest
			Processor1_instruction_master_read                        : in  std_logic                     := 'X';             -- read
			Processor1_instruction_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			Processor2_data_master_address                            : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			Processor2_data_master_waitrequest                        : out std_logic;                                        -- waitrequest
			Processor2_data_master_byteenable                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Processor2_data_master_read                               : in  std_logic                     := 'X';             -- read
			Processor2_data_master_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			Processor2_data_master_write                              : in  std_logic                     := 'X';             -- write
			Processor2_data_master_writedata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Processor2_data_master_debugaccess                        : in  std_logic                     := 'X';             -- debugaccess
			Processor2_instruction_master_address                     : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			Processor2_instruction_master_waitrequest                 : out std_logic;                                        -- waitrequest
			Processor2_instruction_master_read                        : in  std_logic                     := 'X';             -- read
			Processor2_instruction_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			Audio_Subsystem_audio_slave_address                       : out std_logic_vector(1 downto 0);                     -- address
			Audio_Subsystem_audio_slave_write                         : out std_logic;                                        -- write
			Audio_Subsystem_audio_slave_read                          : out std_logic;                                        -- read
			Audio_Subsystem_audio_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Audio_Subsystem_audio_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			Audio_Subsystem_audio_slave_chipselect                    : out std_logic;                                        -- chipselect
			AV_Config_avalon_av_config_slave_address                  : out std_logic_vector(1 downto 0);                     -- address
			AV_Config_avalon_av_config_slave_write                    : out std_logic;                                        -- write
			AV_Config_avalon_av_config_slave_read                     : out std_logic;                                        -- read
			AV_Config_avalon_av_config_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			AV_Config_avalon_av_config_slave_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			AV_Config_avalon_av_config_slave_byteenable               : out std_logic_vector(3 downto 0);                     -- byteenable
			AV_Config_avalon_av_config_slave_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			CameraD5M_0_camera_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Expansion_JP5_avalon_parallel_port_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			Expansion_JP5_avalon_parallel_port_slave_write            : out std_logic;                                        -- write
			Expansion_JP5_avalon_parallel_port_slave_read             : out std_logic;                                        -- read
			Expansion_JP5_avalon_parallel_port_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Expansion_JP5_avalon_parallel_port_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			Expansion_JP5_avalon_parallel_port_slave_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			Expansion_JP5_avalon_parallel_port_slave_chipselect       : out std_logic;                                        -- chipselect
			Flash_flash_data_address                                  : out std_logic_vector(20 downto 0);                    -- address
			Flash_flash_data_write                                    : out std_logic;                                        -- write
			Flash_flash_data_read                                     : out std_logic;                                        -- read
			Flash_flash_data_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Flash_flash_data_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			Flash_flash_data_byteenable                               : out std_logic_vector(3 downto 0);                     -- byteenable
			Flash_flash_data_waitrequest                              : in  std_logic                     := 'X';             -- waitrequest
			Flash_flash_data_chipselect                               : out std_logic;                                        -- chipselect
			Flash_flash_erase_control_write                           : out std_logic;                                        -- write
			Flash_flash_erase_control_read                            : out std_logic;                                        -- read
			Flash_flash_erase_control_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Flash_flash_erase_control_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			Flash_flash_erase_control_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			Flash_flash_erase_control_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			Flash_flash_erase_control_chipselect                      : out std_logic;                                        -- chipselect
			Green_LEDs_avalon_parallel_port_slave_address             : out std_logic_vector(1 downto 0);                     -- address
			Green_LEDs_avalon_parallel_port_slave_write               : out std_logic;                                        -- write
			Green_LEDs_avalon_parallel_port_slave_read                : out std_logic;                                        -- read
			Green_LEDs_avalon_parallel_port_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Green_LEDs_avalon_parallel_port_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			Green_LEDs_avalon_parallel_port_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			Green_LEDs_avalon_parallel_port_slave_chipselect          : out std_logic;                                        -- chipselect
			Interval_Timer_s1_address                                 : out std_logic_vector(2 downto 0);                     -- address
			Interval_Timer_s1_write                                   : out std_logic;                                        -- write
			Interval_Timer_s1_readdata                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Interval_Timer_s1_writedata                               : out std_logic_vector(15 downto 0);                    -- writedata
			Interval_Timer_s1_chipselect                              : out std_logic;                                        -- chipselect
			JTAG_UART_avalon_jtag_slave_address                       : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write                         : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read                          : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect                    : out std_logic;                                        -- chipselect
			JTAG_UART_2nd_Core_avalon_jtag_slave_address              : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_2nd_Core_avalon_jtag_slave_write                : out std_logic;                                        -- write
			JTAG_UART_2nd_Core_avalon_jtag_slave_read                 : out std_logic;                                        -- read
			JTAG_UART_2nd_Core_avalon_jtag_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_2nd_Core_avalon_jtag_slave_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect           : out std_logic;                                        -- chipselect
			Processor1_debug_mem_slave_address                        : out std_logic_vector(8 downto 0);                     -- address
			Processor1_debug_mem_slave_write                          : out std_logic;                                        -- write
			Processor1_debug_mem_slave_read                           : out std_logic;                                        -- read
			Processor1_debug_mem_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Processor1_debug_mem_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			Processor1_debug_mem_slave_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			Processor1_debug_mem_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			Processor1_debug_mem_slave_debugaccess                    : out std_logic;                                        -- debugaccess
			Processor2_debug_mem_slave_address                        : out std_logic_vector(8 downto 0);                     -- address
			Processor2_debug_mem_slave_write                          : out std_logic;                                        -- write
			Processor2_debug_mem_slave_read                           : out std_logic;                                        -- read
			Processor2_debug_mem_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Processor2_debug_mem_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			Processor2_debug_mem_slave_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			Processor2_debug_mem_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			Processor2_debug_mem_slave_debugaccess                    : out std_logic;                                        -- debugaccess
			Pushbuttons_avalon_parallel_port_slave_address            : out std_logic_vector(1 downto 0);                     -- address
			Pushbuttons_avalon_parallel_port_slave_write              : out std_logic;                                        -- write
			Pushbuttons_avalon_parallel_port_slave_read               : out std_logic;                                        -- read
			Pushbuttons_avalon_parallel_port_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Pushbuttons_avalon_parallel_port_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			Pushbuttons_avalon_parallel_port_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			Pushbuttons_avalon_parallel_port_slave_chipselect         : out std_logic;                                        -- chipselect
			Red_LEDs_avalon_parallel_port_slave_address               : out std_logic_vector(1 downto 0);                     -- address
			Red_LEDs_avalon_parallel_port_slave_write                 : out std_logic;                                        -- write
			Red_LEDs_avalon_parallel_port_slave_read                  : out std_logic;                                        -- read
			Red_LEDs_avalon_parallel_port_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Red_LEDs_avalon_parallel_port_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			Red_LEDs_avalon_parallel_port_slave_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			Red_LEDs_avalon_parallel_port_slave_chipselect            : out std_logic;                                        -- chipselect
			SDRAM_s1_address                                          : out std_logic_vector(24 downto 0);                    -- address
			SDRAM_s1_write                                            : out std_logic;                                        -- write
			SDRAM_s1_read                                             : out std_logic;                                        -- read
			SDRAM_s1_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SDRAM_s1_writedata                                        : out std_logic_vector(31 downto 0);                    -- writedata
			SDRAM_s1_byteenable                                       : out std_logic_vector(3 downto 0);                     -- byteenable
			SDRAM_s1_readdatavalid                                    : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                                      : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_s1_chipselect                                       : out std_logic;                                        -- chipselect
			Serial_Port_avalon_rs232_slave_address                    : out std_logic_vector(0 downto 0);                     -- address
			Serial_Port_avalon_rs232_slave_write                      : out std_logic;                                        -- write
			Serial_Port_avalon_rs232_slave_read                       : out std_logic;                                        -- read
			Serial_Port_avalon_rs232_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Serial_Port_avalon_rs232_slave_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			Serial_Port_avalon_rs232_slave_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			Serial_Port_avalon_rs232_slave_chipselect                 : out std_logic;                                        -- chipselect
			Slider_Switches_avalon_parallel_port_slave_address        : out std_logic_vector(1 downto 0);                     -- address
			Slider_Switches_avalon_parallel_port_slave_write          : out std_logic;                                        -- write
			Slider_Switches_avalon_parallel_port_slave_read           : out std_logic;                                        -- read
			Slider_Switches_avalon_parallel_port_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Slider_Switches_avalon_parallel_port_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			Slider_Switches_avalon_parallel_port_slave_byteenable     : out std_logic_vector(3 downto 0);                     -- byteenable
			Slider_Switches_avalon_parallel_port_slave_chipselect     : out std_logic;                                        -- chipselect
			SRAM_avalon_sram_slave_address                            : out std_logic_vector(19 downto 0);                    -- address
			SRAM_avalon_sram_slave_write                              : out std_logic;                                        -- write
			SRAM_avalon_sram_slave_read                               : out std_logic;                                        -- read
			SRAM_avalon_sram_slave_readdata                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SRAM_avalon_sram_slave_writedata                          : out std_logic_vector(15 downto 0);                    -- writedata
			SRAM_avalon_sram_slave_byteenable                         : out std_logic_vector(1 downto 0);                     -- byteenable
			SRAM_avalon_sram_slave_readdatavalid                      : in  std_logic                     := 'X';             -- readdatavalid
			SysID_control_slave_address                               : out std_logic_vector(0 downto 0);                     -- address
			SysID_control_slave_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component nios_system_mm_interconnect_0;

	component nios_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_system_irq_mapper;

	component nios_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_system_rst_controller;

	component nios_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_system_rst_controller_001;

	signal system_pll_sys_clk_clk                                                        : std_logic;                     -- System_PLL:sys_clk_clk -> [AV_Config:clk, Audio_Subsystem:sys_clk_clk, CameraD5M_0:clk_clk, Expansion_JP5:clk, Flash:i_clock, Green_LEDs:clk, Interval_Timer:clk, JTAG_UART:clk, JTAG_UART_2nd_Core:clk, JTAG_to_FPGA_Bridge:clk_clk, Processor1:clk, Processor2:clk, Pushbuttons:clk, Red_LEDs:clk, SDRAM:clk, SRAM:clk, Serial_Port:clk, Slider_Switches:clk, SysID:clock, irq_mapper:clk, irq_mapper_001:clk, mm_interconnect_0:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk]
	signal system_pll_reset_source_reset                                                 : std_logic;                     -- System_PLL:reset_source_reset -> [JTAG_to_FPGA_Bridge:clk_reset_reset, rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in1, system_pll_reset_source_reset:in]
	signal processor1_custom_instruction_master_readra                                   : std_logic;                     -- Processor1:D_ci_readra -> Processor1_custom_instruction_master_translator:ci_slave_readra
	signal processor1_custom_instruction_master_a                                        : std_logic_vector(4 downto 0);  -- Processor1:D_ci_a -> Processor1_custom_instruction_master_translator:ci_slave_a
	signal processor1_custom_instruction_master_b                                        : std_logic_vector(4 downto 0);  -- Processor1:D_ci_b -> Processor1_custom_instruction_master_translator:ci_slave_b
	signal processor1_custom_instruction_master_c                                        : std_logic_vector(4 downto 0);  -- Processor1:D_ci_c -> Processor1_custom_instruction_master_translator:ci_slave_c
	signal processor1_custom_instruction_master_readrb                                   : std_logic;                     -- Processor1:D_ci_readrb -> Processor1_custom_instruction_master_translator:ci_slave_readrb
	signal processor1_custom_instruction_master_clk                                      : std_logic;                     -- Processor1:E_ci_multi_clock -> Processor1_custom_instruction_master_translator:ci_slave_multi_clk
	signal processor1_custom_instruction_master_ipending                                 : std_logic_vector(31 downto 0); -- Processor1:W_ci_ipending -> Processor1_custom_instruction_master_translator:ci_slave_ipending
	signal processor1_custom_instruction_master_start                                    : std_logic;                     -- Processor1:E_ci_multi_start -> Processor1_custom_instruction_master_translator:ci_slave_multi_start
	signal processor1_custom_instruction_master_reset_req                                : std_logic;                     -- Processor1:E_ci_multi_reset_req -> Processor1_custom_instruction_master_translator:ci_slave_multi_reset_req
	signal processor1_custom_instruction_master_done                                     : std_logic;                     -- Processor1_custom_instruction_master_translator:ci_slave_multi_done -> Processor1:E_ci_multi_done
	signal processor1_custom_instruction_master_n                                        : std_logic_vector(7 downto 0);  -- Processor1:D_ci_n -> Processor1_custom_instruction_master_translator:ci_slave_n
	signal processor1_custom_instruction_master_result                                   : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_translator:ci_slave_result -> Processor1:E_ci_result
	signal processor1_custom_instruction_master_estatus                                  : std_logic;                     -- Processor1:W_ci_estatus -> Processor1_custom_instruction_master_translator:ci_slave_estatus
	signal processor1_custom_instruction_master_clk_en                                   : std_logic;                     -- Processor1:E_ci_multi_clk_en -> Processor1_custom_instruction_master_translator:ci_slave_multi_clken
	signal processor1_custom_instruction_master_datab                                    : std_logic_vector(31 downto 0); -- Processor1:E_ci_datab -> Processor1_custom_instruction_master_translator:ci_slave_datab
	signal processor1_custom_instruction_master_dataa                                    : std_logic_vector(31 downto 0); -- Processor1:E_ci_dataa -> Processor1_custom_instruction_master_translator:ci_slave_dataa
	signal processor1_custom_instruction_master_reset                                    : std_logic;                     -- Processor1:E_ci_multi_reset -> Processor1_custom_instruction_master_translator:ci_slave_multi_reset
	signal processor1_custom_instruction_master_writerc                                  : std_logic;                     -- Processor1:D_ci_writerc -> Processor1_custom_instruction_master_translator:ci_slave_writerc
	signal processor1_custom_instruction_master_translator_multi_ci_master_readra        : std_logic;                     -- Processor1_custom_instruction_master_translator:multi_ci_master_readra -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_readra
	signal processor1_custom_instruction_master_translator_multi_ci_master_a             : std_logic_vector(4 downto 0);  -- Processor1_custom_instruction_master_translator:multi_ci_master_a -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_a
	signal processor1_custom_instruction_master_translator_multi_ci_master_b             : std_logic_vector(4 downto 0);  -- Processor1_custom_instruction_master_translator:multi_ci_master_b -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_b
	signal processor1_custom_instruction_master_translator_multi_ci_master_clk           : std_logic;                     -- Processor1_custom_instruction_master_translator:multi_ci_master_clk -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_clk
	signal processor1_custom_instruction_master_translator_multi_ci_master_readrb        : std_logic;                     -- Processor1_custom_instruction_master_translator:multi_ci_master_readrb -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_readrb
	signal processor1_custom_instruction_master_translator_multi_ci_master_c             : std_logic_vector(4 downto 0);  -- Processor1_custom_instruction_master_translator:multi_ci_master_c -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_c
	signal processor1_custom_instruction_master_translator_multi_ci_master_start         : std_logic;                     -- Processor1_custom_instruction_master_translator:multi_ci_master_start -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_start
	signal processor1_custom_instruction_master_translator_multi_ci_master_reset_req     : std_logic;                     -- Processor1_custom_instruction_master_translator:multi_ci_master_reset_req -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	signal processor1_custom_instruction_master_translator_multi_ci_master_done          : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_slave_done -> Processor1_custom_instruction_master_translator:multi_ci_master_done
	signal processor1_custom_instruction_master_translator_multi_ci_master_n             : std_logic_vector(7 downto 0);  -- Processor1_custom_instruction_master_translator:multi_ci_master_n -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_n
	signal processor1_custom_instruction_master_translator_multi_ci_master_result        : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_multi_xconnect:ci_slave_result -> Processor1_custom_instruction_master_translator:multi_ci_master_result
	signal processor1_custom_instruction_master_translator_multi_ci_master_clk_en        : std_logic;                     -- Processor1_custom_instruction_master_translator:multi_ci_master_clken -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_clken
	signal processor1_custom_instruction_master_translator_multi_ci_master_datab         : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_translator:multi_ci_master_datab -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_datab
	signal processor1_custom_instruction_master_translator_multi_ci_master_dataa         : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_translator:multi_ci_master_dataa -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_dataa
	signal processor1_custom_instruction_master_translator_multi_ci_master_reset         : std_logic;                     -- Processor1_custom_instruction_master_translator:multi_ci_master_reset -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_reset
	signal processor1_custom_instruction_master_translator_multi_ci_master_writerc       : std_logic;                     -- Processor1_custom_instruction_master_translator:multi_ci_master_writerc -> Processor1_custom_instruction_master_multi_xconnect:ci_slave_writerc
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_readra         : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_readra -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_a              : std_logic_vector(4 downto 0);  -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_a -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_a
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_b              : std_logic_vector(4 downto 0);  -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_b -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_b
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_readrb         : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_c              : std_logic_vector(4 downto 0);  -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_c -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_c
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_clk            : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_clk -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_ipending       : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_start          : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_start -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_start
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_reset_req      : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_done           : std_logic;                     -- Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Processor1_custom_instruction_master_multi_xconnect:ci_master0_done
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_n              : std_logic_vector(7 downto 0);  -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_n -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_n
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_result         : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Processor1_custom_instruction_master_multi_xconnect:ci_master0_result
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_estatus        : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_clk_en         : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_clken -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_datab          : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_datab -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_dataa          : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_reset          : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_reset -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	signal processor1_custom_instruction_master_multi_xconnect_ci_master0_writerc        : std_logic;                     -- Processor1_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Processor1_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	signal processor1_custom_instruction_master_multi_slave_translator0_ci_master_result : std_logic_vector(31 downto 0); -- Nios2_Floating_Point:result -> Processor1_custom_instruction_master_multi_slave_translator0:ci_master_result
	signal processor1_custom_instruction_master_multi_slave_translator0_ci_master_clk    : std_logic;                     -- Processor1_custom_instruction_master_multi_slave_translator0:ci_master_clk -> Nios2_Floating_Point:clk
	signal processor1_custom_instruction_master_multi_slave_translator0_ci_master_clk_en : std_logic;                     -- Processor1_custom_instruction_master_multi_slave_translator0:ci_master_clken -> Nios2_Floating_Point:clk_en
	signal processor1_custom_instruction_master_multi_slave_translator0_ci_master_datab  : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_multi_slave_translator0:ci_master_datab -> Nios2_Floating_Point:datab
	signal processor1_custom_instruction_master_multi_slave_translator0_ci_master_dataa  : std_logic_vector(31 downto 0); -- Processor1_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> Nios2_Floating_Point:dataa
	signal processor1_custom_instruction_master_multi_slave_translator0_ci_master_start  : std_logic;                     -- Processor1_custom_instruction_master_multi_slave_translator0:ci_master_start -> Nios2_Floating_Point:start
	signal processor1_custom_instruction_master_multi_slave_translator0_ci_master_reset  : std_logic;                     -- Processor1_custom_instruction_master_multi_slave_translator0:ci_master_reset -> Nios2_Floating_Point:reset
	signal processor1_custom_instruction_master_multi_slave_translator0_ci_master_done   : std_logic;                     -- Nios2_Floating_Point:done -> Processor1_custom_instruction_master_multi_slave_translator0:ci_master_done
	signal processor1_custom_instruction_master_multi_slave_translator0_ci_master_n      : std_logic_vector(1 downto 0);  -- Processor1_custom_instruction_master_multi_slave_translator0:ci_master_n -> Nios2_Floating_Point:n
	signal processor2_custom_instruction_master_readra                                   : std_logic;                     -- Processor2:D_ci_readra -> Processor2_custom_instruction_master_translator:ci_slave_readra
	signal processor2_custom_instruction_master_a                                        : std_logic_vector(4 downto 0);  -- Processor2:D_ci_a -> Processor2_custom_instruction_master_translator:ci_slave_a
	signal processor2_custom_instruction_master_b                                        : std_logic_vector(4 downto 0);  -- Processor2:D_ci_b -> Processor2_custom_instruction_master_translator:ci_slave_b
	signal processor2_custom_instruction_master_c                                        : std_logic_vector(4 downto 0);  -- Processor2:D_ci_c -> Processor2_custom_instruction_master_translator:ci_slave_c
	signal processor2_custom_instruction_master_readrb                                   : std_logic;                     -- Processor2:D_ci_readrb -> Processor2_custom_instruction_master_translator:ci_slave_readrb
	signal processor2_custom_instruction_master_clk                                      : std_logic;                     -- Processor2:E_ci_multi_clock -> Processor2_custom_instruction_master_translator:ci_slave_multi_clk
	signal processor2_custom_instruction_master_ipending                                 : std_logic_vector(31 downto 0); -- Processor2:W_ci_ipending -> Processor2_custom_instruction_master_translator:ci_slave_ipending
	signal processor2_custom_instruction_master_start                                    : std_logic;                     -- Processor2:E_ci_multi_start -> Processor2_custom_instruction_master_translator:ci_slave_multi_start
	signal processor2_custom_instruction_master_reset_req                                : std_logic;                     -- Processor2:E_ci_multi_reset_req -> Processor2_custom_instruction_master_translator:ci_slave_multi_reset_req
	signal processor2_custom_instruction_master_done                                     : std_logic;                     -- Processor2_custom_instruction_master_translator:ci_slave_multi_done -> Processor2:E_ci_multi_done
	signal processor2_custom_instruction_master_n                                        : std_logic_vector(7 downto 0);  -- Processor2:D_ci_n -> Processor2_custom_instruction_master_translator:ci_slave_n
	signal processor2_custom_instruction_master_result                                   : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_translator:ci_slave_result -> Processor2:E_ci_result
	signal processor2_custom_instruction_master_estatus                                  : std_logic;                     -- Processor2:W_ci_estatus -> Processor2_custom_instruction_master_translator:ci_slave_estatus
	signal processor2_custom_instruction_master_clk_en                                   : std_logic;                     -- Processor2:E_ci_multi_clk_en -> Processor2_custom_instruction_master_translator:ci_slave_multi_clken
	signal processor2_custom_instruction_master_datab                                    : std_logic_vector(31 downto 0); -- Processor2:E_ci_datab -> Processor2_custom_instruction_master_translator:ci_slave_datab
	signal processor2_custom_instruction_master_dataa                                    : std_logic_vector(31 downto 0); -- Processor2:E_ci_dataa -> Processor2_custom_instruction_master_translator:ci_slave_dataa
	signal processor2_custom_instruction_master_reset                                    : std_logic;                     -- Processor2:E_ci_multi_reset -> Processor2_custom_instruction_master_translator:ci_slave_multi_reset
	signal processor2_custom_instruction_master_writerc                                  : std_logic;                     -- Processor2:D_ci_writerc -> Processor2_custom_instruction_master_translator:ci_slave_writerc
	signal processor2_custom_instruction_master_translator_multi_ci_master_readra        : std_logic;                     -- Processor2_custom_instruction_master_translator:multi_ci_master_readra -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_readra
	signal processor2_custom_instruction_master_translator_multi_ci_master_a             : std_logic_vector(4 downto 0);  -- Processor2_custom_instruction_master_translator:multi_ci_master_a -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_a
	signal processor2_custom_instruction_master_translator_multi_ci_master_b             : std_logic_vector(4 downto 0);  -- Processor2_custom_instruction_master_translator:multi_ci_master_b -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_b
	signal processor2_custom_instruction_master_translator_multi_ci_master_clk           : std_logic;                     -- Processor2_custom_instruction_master_translator:multi_ci_master_clk -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_clk
	signal processor2_custom_instruction_master_translator_multi_ci_master_readrb        : std_logic;                     -- Processor2_custom_instruction_master_translator:multi_ci_master_readrb -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_readrb
	signal processor2_custom_instruction_master_translator_multi_ci_master_c             : std_logic_vector(4 downto 0);  -- Processor2_custom_instruction_master_translator:multi_ci_master_c -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_c
	signal processor2_custom_instruction_master_translator_multi_ci_master_start         : std_logic;                     -- Processor2_custom_instruction_master_translator:multi_ci_master_start -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_start
	signal processor2_custom_instruction_master_translator_multi_ci_master_reset_req     : std_logic;                     -- Processor2_custom_instruction_master_translator:multi_ci_master_reset_req -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	signal processor2_custom_instruction_master_translator_multi_ci_master_done          : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_slave_done -> Processor2_custom_instruction_master_translator:multi_ci_master_done
	signal processor2_custom_instruction_master_translator_multi_ci_master_n             : std_logic_vector(7 downto 0);  -- Processor2_custom_instruction_master_translator:multi_ci_master_n -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_n
	signal processor2_custom_instruction_master_translator_multi_ci_master_result        : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_multi_xconnect:ci_slave_result -> Processor2_custom_instruction_master_translator:multi_ci_master_result
	signal processor2_custom_instruction_master_translator_multi_ci_master_clk_en        : std_logic;                     -- Processor2_custom_instruction_master_translator:multi_ci_master_clken -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_clken
	signal processor2_custom_instruction_master_translator_multi_ci_master_datab         : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_translator:multi_ci_master_datab -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_datab
	signal processor2_custom_instruction_master_translator_multi_ci_master_dataa         : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_translator:multi_ci_master_dataa -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_dataa
	signal processor2_custom_instruction_master_translator_multi_ci_master_reset         : std_logic;                     -- Processor2_custom_instruction_master_translator:multi_ci_master_reset -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_reset
	signal processor2_custom_instruction_master_translator_multi_ci_master_writerc       : std_logic;                     -- Processor2_custom_instruction_master_translator:multi_ci_master_writerc -> Processor2_custom_instruction_master_multi_xconnect:ci_slave_writerc
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_readra         : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_readra -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_a              : std_logic_vector(4 downto 0);  -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_a -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_a
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_b              : std_logic_vector(4 downto 0);  -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_b -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_b
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_readrb         : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_c              : std_logic_vector(4 downto 0);  -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_c -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_c
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_clk            : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_clk -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_ipending       : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_start          : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_start -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_start
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_reset_req      : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_done           : std_logic;                     -- Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Processor2_custom_instruction_master_multi_xconnect:ci_master0_done
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_n              : std_logic_vector(7 downto 0);  -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_n -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_n
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_result         : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Processor2_custom_instruction_master_multi_xconnect:ci_master0_result
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_estatus        : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_clk_en         : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_clken -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_datab          : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_datab -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_dataa          : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_reset          : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_reset -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	signal processor2_custom_instruction_master_multi_xconnect_ci_master0_writerc        : std_logic;                     -- Processor2_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Processor2_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	signal processor2_custom_instruction_master_multi_slave_translator0_ci_master_result : std_logic_vector(31 downto 0); -- Nios2_Floating_Point_2nd_Core:result -> Processor2_custom_instruction_master_multi_slave_translator0:ci_master_result
	signal processor2_custom_instruction_master_multi_slave_translator0_ci_master_clk    : std_logic;                     -- Processor2_custom_instruction_master_multi_slave_translator0:ci_master_clk -> Nios2_Floating_Point_2nd_Core:clk
	signal processor2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en : std_logic;                     -- Processor2_custom_instruction_master_multi_slave_translator0:ci_master_clken -> Nios2_Floating_Point_2nd_Core:clk_en
	signal processor2_custom_instruction_master_multi_slave_translator0_ci_master_datab  : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_multi_slave_translator0:ci_master_datab -> Nios2_Floating_Point_2nd_Core:datab
	signal processor2_custom_instruction_master_multi_slave_translator0_ci_master_dataa  : std_logic_vector(31 downto 0); -- Processor2_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> Nios2_Floating_Point_2nd_Core:dataa
	signal processor2_custom_instruction_master_multi_slave_translator0_ci_master_start  : std_logic;                     -- Processor2_custom_instruction_master_multi_slave_translator0:ci_master_start -> Nios2_Floating_Point_2nd_Core:start
	signal processor2_custom_instruction_master_multi_slave_translator0_ci_master_reset  : std_logic;                     -- Processor2_custom_instruction_master_multi_slave_translator0:ci_master_reset -> Nios2_Floating_Point_2nd_Core:reset
	signal processor2_custom_instruction_master_multi_slave_translator0_ci_master_done   : std_logic;                     -- Nios2_Floating_Point_2nd_Core:done -> Processor2_custom_instruction_master_multi_slave_translator0:ci_master_done
	signal processor2_custom_instruction_master_multi_slave_translator0_ci_master_n      : std_logic_vector(1 downto 0);  -- Processor2_custom_instruction_master_multi_slave_translator0:ci_master_n -> Nios2_Floating_Point_2nd_Core:n
	signal processor2_data_master_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor2_data_master_readdata -> Processor2:d_readdata
	signal processor2_data_master_waitrequest                                            : std_logic;                     -- mm_interconnect_0:Processor2_data_master_waitrequest -> Processor2:d_waitrequest
	signal processor2_data_master_debugaccess                                            : std_logic;                     -- Processor2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Processor2_data_master_debugaccess
	signal processor2_data_master_address                                                : std_logic_vector(28 downto 0); -- Processor2:d_address -> mm_interconnect_0:Processor2_data_master_address
	signal processor2_data_master_byteenable                                             : std_logic_vector(3 downto 0);  -- Processor2:d_byteenable -> mm_interconnect_0:Processor2_data_master_byteenable
	signal processor2_data_master_read                                                   : std_logic;                     -- Processor2:d_read -> mm_interconnect_0:Processor2_data_master_read
	signal processor2_data_master_write                                                  : std_logic;                     -- Processor2:d_write -> mm_interconnect_0:Processor2_data_master_write
	signal processor2_data_master_writedata                                              : std_logic_vector(31 downto 0); -- Processor2:d_writedata -> mm_interconnect_0:Processor2_data_master_writedata
	signal processor1_data_master_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor1_data_master_readdata -> Processor1:d_readdata
	signal processor1_data_master_waitrequest                                            : std_logic;                     -- mm_interconnect_0:Processor1_data_master_waitrequest -> Processor1:d_waitrequest
	signal processor1_data_master_debugaccess                                            : std_logic;                     -- Processor1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Processor1_data_master_debugaccess
	signal processor1_data_master_address                                                : std_logic_vector(28 downto 0); -- Processor1:d_address -> mm_interconnect_0:Processor1_data_master_address
	signal processor1_data_master_byteenable                                             : std_logic_vector(3 downto 0);  -- Processor1:d_byteenable -> mm_interconnect_0:Processor1_data_master_byteenable
	signal processor1_data_master_read                                                   : std_logic;                     -- Processor1:d_read -> mm_interconnect_0:Processor1_data_master_read
	signal processor1_data_master_write                                                  : std_logic;                     -- Processor1:d_write -> mm_interconnect_0:Processor1_data_master_write
	signal processor1_data_master_writedata                                              : std_logic_vector(31 downto 0); -- Processor1:d_writedata -> mm_interconnect_0:Processor1_data_master_writedata
	signal jtag_to_fpga_bridge_master_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdata -> JTAG_to_FPGA_Bridge:master_readdata
	signal jtag_to_fpga_bridge_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:JTAG_to_FPGA_Bridge_master_waitrequest -> JTAG_to_FPGA_Bridge:master_waitrequest
	signal jtag_to_fpga_bridge_master_address                                            : std_logic_vector(31 downto 0); -- JTAG_to_FPGA_Bridge:master_address -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_address
	signal jtag_to_fpga_bridge_master_read                                               : std_logic;                     -- JTAG_to_FPGA_Bridge:master_read -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_read
	signal jtag_to_fpga_bridge_master_byteenable                                         : std_logic_vector(3 downto 0);  -- JTAG_to_FPGA_Bridge:master_byteenable -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_byteenable
	signal jtag_to_fpga_bridge_master_readdatavalid                                      : std_logic;                     -- mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdatavalid -> JTAG_to_FPGA_Bridge:master_readdatavalid
	signal jtag_to_fpga_bridge_master_write                                              : std_logic;                     -- JTAG_to_FPGA_Bridge:master_write -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_write
	signal jtag_to_fpga_bridge_master_writedata                                          : std_logic_vector(31 downto 0); -- JTAG_to_FPGA_Bridge:master_writedata -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_writedata
	signal processor1_instruction_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor1_instruction_master_readdata -> Processor1:i_readdata
	signal processor1_instruction_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:Processor1_instruction_master_waitrequest -> Processor1:i_waitrequest
	signal processor1_instruction_master_address                                         : std_logic_vector(27 downto 0); -- Processor1:i_address -> mm_interconnect_0:Processor1_instruction_master_address
	signal processor1_instruction_master_read                                            : std_logic;                     -- Processor1:i_read -> mm_interconnect_0:Processor1_instruction_master_read
	signal processor2_instruction_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor2_instruction_master_readdata -> Processor2:i_readdata
	signal processor2_instruction_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:Processor2_instruction_master_waitrequest -> Processor2:i_waitrequest
	signal processor2_instruction_master_address                                         : std_logic_vector(27 downto 0); -- Processor2:i_address -> mm_interconnect_0:Processor2_instruction_master_address
	signal processor2_instruction_master_read                                            : std_logic;                     -- Processor2:i_read -> mm_interconnect_0:Processor2_instruction_master_read
	signal mm_interconnect_0_audio_subsystem_audio_slave_chipselect                      : std_logic;                     -- mm_interconnect_0:Audio_Subsystem_audio_slave_chipselect -> Audio_Subsystem:audio_slave_chipselect
	signal mm_interconnect_0_audio_subsystem_audio_slave_readdata                        : std_logic_vector(31 downto 0); -- Audio_Subsystem:audio_slave_readdata -> mm_interconnect_0:Audio_Subsystem_audio_slave_readdata
	signal mm_interconnect_0_audio_subsystem_audio_slave_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Audio_Subsystem_audio_slave_address -> Audio_Subsystem:audio_slave_address
	signal mm_interconnect_0_audio_subsystem_audio_slave_read                            : std_logic;                     -- mm_interconnect_0:Audio_Subsystem_audio_slave_read -> Audio_Subsystem:audio_slave_read
	signal mm_interconnect_0_audio_subsystem_audio_slave_write                           : std_logic;                     -- mm_interconnect_0:Audio_Subsystem_audio_slave_write -> Audio_Subsystem:audio_slave_write
	signal mm_interconnect_0_audio_subsystem_audio_slave_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Audio_Subsystem_audio_slave_writedata -> Audio_Subsystem:audio_slave_writedata
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect             : std_logic;                     -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect -> JTAG_UART_2nd_Core:av_chipselect
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata               : std_logic_vector(31 downto 0); -- JTAG_UART_2nd_Core:av_readdata -> mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest            : std_logic;                     -- JTAG_UART_2nd_Core:av_waitrequest -> mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_address -> JTAG_UART_2nd_Core:av_address
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read                   : std_logic;                     -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write                  : std_logic;                     -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_writedata -> JTAG_UART_2nd_Core:av_writedata
	signal mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_chipselect         : std_logic;                     -- mm_interconnect_0:Expansion_JP5_avalon_parallel_port_slave_chipselect -> Expansion_JP5:chipselect
	signal mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_readdata           : std_logic_vector(31 downto 0); -- Expansion_JP5:readdata -> mm_interconnect_0:Expansion_JP5_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Expansion_JP5_avalon_parallel_port_slave_address -> Expansion_JP5:address
	signal mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_read               : std_logic;                     -- mm_interconnect_0:Expansion_JP5_avalon_parallel_port_slave_read -> Expansion_JP5:read
	signal mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Expansion_JP5_avalon_parallel_port_slave_byteenable -> Expansion_JP5:byteenable
	signal mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_write              : std_logic;                     -- mm_interconnect_0:Expansion_JP5_avalon_parallel_port_slave_write -> Expansion_JP5:write
	signal mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:Expansion_JP5_avalon_parallel_port_slave_writedata -> Expansion_JP5:writedata
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect           : std_logic;                     -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_chipselect -> Pushbuttons:chipselect
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata             : std_logic_vector(31 downto 0); -- Pushbuttons:readdata -> mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_address -> Pushbuttons:address
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read                 : std_logic;                     -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_read -> Pushbuttons:read
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_byteenable -> Pushbuttons:byteenable
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write                : std_logic;                     -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_write -> Pushbuttons:write
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_writedata -> Pushbuttons:writedata
	signal mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect                   : std_logic;                     -- mm_interconnect_0:Serial_Port_avalon_rs232_slave_chipselect -> Serial_Port:chipselect
	signal mm_interconnect_0_serial_port_avalon_rs232_slave_readdata                     : std_logic_vector(31 downto 0); -- Serial_Port:readdata -> mm_interconnect_0:Serial_Port_avalon_rs232_slave_readdata
	signal mm_interconnect_0_serial_port_avalon_rs232_slave_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:Serial_Port_avalon_rs232_slave_address -> Serial_Port:address
	signal mm_interconnect_0_serial_port_avalon_rs232_slave_read                         : std_logic;                     -- mm_interconnect_0:Serial_Port_avalon_rs232_slave_read -> Serial_Port:read
	signal mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Serial_Port_avalon_rs232_slave_byteenable -> Serial_Port:byteenable
	signal mm_interconnect_0_serial_port_avalon_rs232_slave_write                        : std_logic;                     -- mm_interconnect_0:Serial_Port_avalon_rs232_slave_write -> Serial_Port:write
	signal mm_interconnect_0_serial_port_avalon_rs232_slave_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:Serial_Port_avalon_rs232_slave_writedata -> Serial_Port:writedata
	signal mm_interconnect_0_camerad5m_0_camera_slave_readdata                           : std_logic_vector(31 downto 0); -- CameraD5M_0:camera_slave_readdata -> mm_interconnect_0:CameraD5M_0_camera_slave_readdata
	signal mm_interconnect_0_processor2_debug_mem_slave_readdata                         : std_logic_vector(31 downto 0); -- Processor2:debug_mem_slave_readdata -> mm_interconnect_0:Processor2_debug_mem_slave_readdata
	signal mm_interconnect_0_processor2_debug_mem_slave_waitrequest                      : std_logic;                     -- Processor2:debug_mem_slave_waitrequest -> mm_interconnect_0:Processor2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_processor2_debug_mem_slave_debugaccess                      : std_logic;                     -- mm_interconnect_0:Processor2_debug_mem_slave_debugaccess -> Processor2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_processor2_debug_mem_slave_address                          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Processor2_debug_mem_slave_address -> Processor2:debug_mem_slave_address
	signal mm_interconnect_0_processor2_debug_mem_slave_read                             : std_logic;                     -- mm_interconnect_0:Processor2_debug_mem_slave_read -> Processor2:debug_mem_slave_read
	signal mm_interconnect_0_processor2_debug_mem_slave_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Processor2_debug_mem_slave_byteenable -> Processor2:debug_mem_slave_byteenable
	signal mm_interconnect_0_processor2_debug_mem_slave_write                            : std_logic;                     -- mm_interconnect_0:Processor2_debug_mem_slave_write -> Processor2:debug_mem_slave_write
	signal mm_interconnect_0_processor2_debug_mem_slave_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor2_debug_mem_slave_writedata -> Processor2:debug_mem_slave_writedata
	signal mm_interconnect_0_interval_timer_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:Interval_Timer_s1_chipselect -> Interval_Timer:chipselect
	signal mm_interconnect_0_interval_timer_s1_readdata                                  : std_logic_vector(15 downto 0); -- Interval_Timer:readdata -> mm_interconnect_0:Interval_Timer_s1_readdata
	signal mm_interconnect_0_interval_timer_s1_address                                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Interval_Timer_s1_address -> Interval_Timer:address
	signal mm_interconnect_0_interval_timer_s1_write                                     : std_logic;                     -- mm_interconnect_0:Interval_Timer_s1_write -> mm_interconnect_0_interval_timer_s1_write:in
	signal mm_interconnect_0_interval_timer_s1_writedata                                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:Interval_Timer_s1_writedata -> Interval_Timer:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                                         : std_logic;                     -- mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                           : std_logic_vector(31 downto 0); -- SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                        : std_logic;                     -- SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                            : std_logic_vector(24 downto 0); -- mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_0_sdram_s1_read                                               : std_logic;                     -- mm_interconnect_0:SDRAM_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SDRAM_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                                      : std_logic;                     -- SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                              : std_logic;                     -- mm_interconnect_0:SDRAM_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	signal mm_interconnect_0_av_config_avalon_av_config_slave_readdata                   : std_logic_vector(31 downto 0); -- AV_Config:readdata -> mm_interconnect_0:AV_Config_avalon_av_config_slave_readdata
	signal mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest                : std_logic;                     -- AV_Config:waitrequest -> mm_interconnect_0:AV_Config_avalon_av_config_slave_waitrequest
	signal mm_interconnect_0_av_config_avalon_av_config_slave_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:AV_Config_avalon_av_config_slave_address -> AV_Config:address
	signal mm_interconnect_0_av_config_avalon_av_config_slave_read                       : std_logic;                     -- mm_interconnect_0:AV_Config_avalon_av_config_slave_read -> AV_Config:read
	signal mm_interconnect_0_av_config_avalon_av_config_slave_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:AV_Config_avalon_av_config_slave_byteenable -> AV_Config:byteenable
	signal mm_interconnect_0_av_config_avalon_av_config_slave_write                      : std_logic;                     -- mm_interconnect_0:AV_Config_avalon_av_config_slave_write -> AV_Config:write
	signal mm_interconnect_0_av_config_avalon_av_config_slave_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:AV_Config_avalon_av_config_slave_writedata -> AV_Config:writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect                      : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                        : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest                     : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                            : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                           : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal mm_interconnect_0_red_leds_avalon_parallel_port_slave_chipselect              : std_logic;                     -- mm_interconnect_0:Red_LEDs_avalon_parallel_port_slave_chipselect -> Red_LEDs:chipselect
	signal mm_interconnect_0_red_leds_avalon_parallel_port_slave_readdata                : std_logic_vector(31 downto 0); -- Red_LEDs:readdata -> mm_interconnect_0:Red_LEDs_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_red_leds_avalon_parallel_port_slave_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Red_LEDs_avalon_parallel_port_slave_address -> Red_LEDs:address
	signal mm_interconnect_0_red_leds_avalon_parallel_port_slave_read                    : std_logic;                     -- mm_interconnect_0:Red_LEDs_avalon_parallel_port_slave_read -> Red_LEDs:read
	signal mm_interconnect_0_red_leds_avalon_parallel_port_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Red_LEDs_avalon_parallel_port_slave_byteenable -> Red_LEDs:byteenable
	signal mm_interconnect_0_red_leds_avalon_parallel_port_slave_write                   : std_logic;                     -- mm_interconnect_0:Red_LEDs_avalon_parallel_port_slave_write -> Red_LEDs:write
	signal mm_interconnect_0_red_leds_avalon_parallel_port_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:Red_LEDs_avalon_parallel_port_slave_writedata -> Red_LEDs:writedata
	signal mm_interconnect_0_green_leds_avalon_parallel_port_slave_chipselect            : std_logic;                     -- mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_chipselect -> Green_LEDs:chipselect
	signal mm_interconnect_0_green_leds_avalon_parallel_port_slave_readdata              : std_logic_vector(31 downto 0); -- Green_LEDs:readdata -> mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_green_leds_avalon_parallel_port_slave_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_address -> Green_LEDs:address
	signal mm_interconnect_0_green_leds_avalon_parallel_port_slave_read                  : std_logic;                     -- mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_read -> Green_LEDs:read
	signal mm_interconnect_0_green_leds_avalon_parallel_port_slave_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_byteenable -> Green_LEDs:byteenable
	signal mm_interconnect_0_green_leds_avalon_parallel_port_slave_write                 : std_logic;                     -- mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_write -> Green_LEDs:write
	signal mm_interconnect_0_green_leds_avalon_parallel_port_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_writedata -> Green_LEDs:writedata
	signal mm_interconnect_0_slider_switches_avalon_parallel_port_slave_chipselect       : std_logic;                     -- mm_interconnect_0:Slider_Switches_avalon_parallel_port_slave_chipselect -> Slider_Switches:chipselect
	signal mm_interconnect_0_slider_switches_avalon_parallel_port_slave_readdata         : std_logic_vector(31 downto 0); -- Slider_Switches:readdata -> mm_interconnect_0:Slider_Switches_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_slider_switches_avalon_parallel_port_slave_address          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Slider_Switches_avalon_parallel_port_slave_address -> Slider_Switches:address
	signal mm_interconnect_0_slider_switches_avalon_parallel_port_slave_read             : std_logic;                     -- mm_interconnect_0:Slider_Switches_avalon_parallel_port_slave_read -> Slider_Switches:read
	signal mm_interconnect_0_slider_switches_avalon_parallel_port_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Slider_Switches_avalon_parallel_port_slave_byteenable -> Slider_Switches:byteenable
	signal mm_interconnect_0_slider_switches_avalon_parallel_port_slave_write            : std_logic;                     -- mm_interconnect_0:Slider_Switches_avalon_parallel_port_slave_write -> Slider_Switches:write
	signal mm_interconnect_0_slider_switches_avalon_parallel_port_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Slider_Switches_avalon_parallel_port_slave_writedata -> Slider_Switches:writedata
	signal mm_interconnect_0_sram_avalon_sram_slave_readdata                             : std_logic_vector(15 downto 0); -- SRAM:readdata -> mm_interconnect_0:SRAM_avalon_sram_slave_readdata
	signal mm_interconnect_0_sram_avalon_sram_slave_address                              : std_logic_vector(19 downto 0); -- mm_interconnect_0:SRAM_avalon_sram_slave_address -> SRAM:address
	signal mm_interconnect_0_sram_avalon_sram_slave_read                                 : std_logic;                     -- mm_interconnect_0:SRAM_avalon_sram_slave_read -> SRAM:read
	signal mm_interconnect_0_sram_avalon_sram_slave_byteenable                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SRAM_avalon_sram_slave_byteenable -> SRAM:byteenable
	signal mm_interconnect_0_sram_avalon_sram_slave_readdatavalid                        : std_logic;                     -- SRAM:readdatavalid -> mm_interconnect_0:SRAM_avalon_sram_slave_readdatavalid
	signal mm_interconnect_0_sram_avalon_sram_slave_write                                : std_logic;                     -- mm_interconnect_0:SRAM_avalon_sram_slave_write -> SRAM:write
	signal mm_interconnect_0_sram_avalon_sram_slave_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:SRAM_avalon_sram_slave_writedata -> SRAM:writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                                : std_logic_vector(31 downto 0); -- SysID:readdata -> mm_interconnect_0:SysID_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:SysID_control_slave_address -> SysID:address
	signal mm_interconnect_0_flash_flash_data_chipselect                                 : std_logic;                     -- mm_interconnect_0:Flash_flash_data_chipselect -> Flash:i_avalon_chip_select
	signal mm_interconnect_0_flash_flash_data_readdata                                   : std_logic_vector(31 downto 0); -- Flash:o_avalon_readdata -> mm_interconnect_0:Flash_flash_data_readdata
	signal mm_interconnect_0_flash_flash_data_waitrequest                                : std_logic;                     -- Flash:o_avalon_waitrequest -> mm_interconnect_0:Flash_flash_data_waitrequest
	signal mm_interconnect_0_flash_flash_data_address                                    : std_logic_vector(20 downto 0); -- mm_interconnect_0:Flash_flash_data_address -> Flash:i_avalon_address
	signal mm_interconnect_0_flash_flash_data_read                                       : std_logic;                     -- mm_interconnect_0:Flash_flash_data_read -> Flash:i_avalon_read
	signal mm_interconnect_0_flash_flash_data_byteenable                                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Flash_flash_data_byteenable -> Flash:i_avalon_byteenable
	signal mm_interconnect_0_flash_flash_data_write                                      : std_logic;                     -- mm_interconnect_0:Flash_flash_data_write -> Flash:i_avalon_write
	signal mm_interconnect_0_flash_flash_data_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:Flash_flash_data_writedata -> Flash:i_avalon_writedata
	signal mm_interconnect_0_flash_flash_erase_control_chipselect                        : std_logic;                     -- mm_interconnect_0:Flash_flash_erase_control_chipselect -> Flash:i_avalon_erase_chip_select
	signal mm_interconnect_0_flash_flash_erase_control_readdata                          : std_logic_vector(31 downto 0); -- Flash:o_avalon_erase_readdata -> mm_interconnect_0:Flash_flash_erase_control_readdata
	signal mm_interconnect_0_flash_flash_erase_control_waitrequest                       : std_logic;                     -- Flash:o_avalon_erase_waitrequest -> mm_interconnect_0:Flash_flash_erase_control_waitrequest
	signal mm_interconnect_0_flash_flash_erase_control_read                              : std_logic;                     -- mm_interconnect_0:Flash_flash_erase_control_read -> Flash:i_avalon_erase_read
	signal mm_interconnect_0_flash_flash_erase_control_byteenable                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Flash_flash_erase_control_byteenable -> Flash:i_avalon_erase_byteenable
	signal mm_interconnect_0_flash_flash_erase_control_write                             : std_logic;                     -- mm_interconnect_0:Flash_flash_erase_control_write -> Flash:i_avalon_erase_write
	signal mm_interconnect_0_flash_flash_erase_control_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:Flash_flash_erase_control_writedata -> Flash:i_avalon_erase_writedata
	signal mm_interconnect_0_processor1_debug_mem_slave_readdata                         : std_logic_vector(31 downto 0); -- Processor1:debug_mem_slave_readdata -> mm_interconnect_0:Processor1_debug_mem_slave_readdata
	signal mm_interconnect_0_processor1_debug_mem_slave_waitrequest                      : std_logic;                     -- Processor1:debug_mem_slave_waitrequest -> mm_interconnect_0:Processor1_debug_mem_slave_waitrequest
	signal mm_interconnect_0_processor1_debug_mem_slave_debugaccess                      : std_logic;                     -- mm_interconnect_0:Processor1_debug_mem_slave_debugaccess -> Processor1:debug_mem_slave_debugaccess
	signal mm_interconnect_0_processor1_debug_mem_slave_address                          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Processor1_debug_mem_slave_address -> Processor1:debug_mem_slave_address
	signal mm_interconnect_0_processor1_debug_mem_slave_read                             : std_logic;                     -- mm_interconnect_0:Processor1_debug_mem_slave_read -> Processor1:debug_mem_slave_read
	signal mm_interconnect_0_processor1_debug_mem_slave_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Processor1_debug_mem_slave_byteenable -> Processor1:debug_mem_slave_byteenable
	signal mm_interconnect_0_processor1_debug_mem_slave_write                            : std_logic;                     -- mm_interconnect_0:Processor1_debug_mem_slave_write -> Processor1:debug_mem_slave_write
	signal mm_interconnect_0_processor1_debug_mem_slave_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor1_debug_mem_slave_writedata -> Processor1:debug_mem_slave_writedata
	signal irq_mapper_receiver5_irq                                                      : std_logic;                     -- JTAG_UART:av_irq -> irq_mapper:receiver5_irq
	signal processor1_irq_irq                                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> Processor1:irq
	signal irq_mapper_001_receiver5_irq                                                  : std_logic;                     -- JTAG_UART_2nd_Core:av_irq -> irq_mapper_001:receiver5_irq
	signal processor2_irq_irq                                                            : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> Processor2:irq
	signal irq_mapper_receiver0_irq                                                      : std_logic;                     -- Audio_Subsystem:audio_irq_irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	signal irq_mapper_receiver1_irq                                                      : std_logic;                     -- Expansion_JP5:irq -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	signal irq_mapper_receiver4_irq                                                      : std_logic;                     -- Interval_Timer:irq -> [irq_mapper:receiver4_irq, irq_mapper_001:receiver4_irq]
	signal irq_mapper_receiver2_irq                                                      : std_logic;                     -- Pushbuttons:irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver2_irq]
	signal irq_mapper_receiver3_irq                                                      : std_logic;                     -- Serial_Port:irq -> [irq_mapper:receiver3_irq, irq_mapper_001:receiver3_irq]
	signal rst_controller_reset_out_reset                                                : std_logic;                     -- rst_controller:reset_out -> [AV_Config:reset, Expansion_JP5:reset, Green_LEDs:reset, Pushbuttons:reset, Red_LEDs:reset, SRAM:reset, Serial_Port:reset, Slider_Switches:reset, mm_interconnect_0:JTAG_UART_2nd_Core_reset_reset_bridge_in_reset_reset, mm_interconnect_0:JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                                            : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:Processor1_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset_req                                        : std_logic;                     -- rst_controller_001:reset_req -> [Processor1:reset_req, rst_translator:reset_req_in]
	signal processor1_debug_reset_request_reset                                          : std_logic;                     -- Processor1:debug_reset_request -> rst_controller_001:reset_in0
	signal rst_controller_002_reset_out_reset                                            : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper_001:reset, mm_interconnect_0:Processor2_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset_req                                        : std_logic;                     -- rst_controller_002:reset_req -> [Processor2:reset_req, rst_translator_001:reset_req_in]
	signal processor2_debug_reset_request_reset                                          : std_logic;                     -- Processor2:debug_reset_request -> rst_controller_002:reset_in0
	signal system_pll_reset_source_reset_ports_inv                                       : std_logic;                     -- system_pll_reset_source_reset:inv -> [Audio_Subsystem:sys_reset_reset_n, CameraD5M_0:reset_reset_n]
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read_ports_inv         : std_logic;                     -- mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read:inv -> JTAG_UART_2nd_Core:av_read_n
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write_ports_inv        : std_logic;                     -- mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write:inv -> JTAG_UART_2nd_Core:av_write_n
	signal mm_interconnect_0_interval_timer_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_interval_timer_s1_write:inv -> Interval_Timer:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                                     : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                               : std_logic_vector(3 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                                    : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv                  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Flash:i_reset_n, Interval_Timer:reset_n, JTAG_UART:rst_n, JTAG_UART_2nd_Core:rst_n, SDRAM:reset_n, SysID:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> Processor1:reset_n
	signal rst_controller_002_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> Processor2:reset_n

begin

	av_config : component nios_system_AV_Config
		port map (
			clk         => system_pll_sys_clk_clk,                                         --                    clk.clk
			reset       => rst_controller_reset_out_reset,                                 --                  reset.reset
			address     => mm_interconnect_0_av_config_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_0_av_config_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_0_av_config_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_0_av_config_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_0_av_config_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_0_av_config_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => av_config_SDAT,                                                 --     external_interface.export
			I2C_SCLK    => av_config_SCLK                                                  --                       .export
		);

	audio_subsystem : component nios_system_Audio_Subsystem
		port map (
			audio_ADCDAT              => audio_ADCDAT,                                             --               audio.ADCDAT
			audio_ADCLRCK             => audio_ADCLRCK,                                            --                    .ADCLRCK
			audio_BCLK                => audio_BCLK,                                               --                    .BCLK
			audio_DACDAT              => audio_DACDAT,                                             --                    .DACDAT
			audio_DACLRCK             => audio_DACLRCK,                                            --                    .DACLRCK
			audio_clk_clk             => audio_clk_clk,                                            --           audio_clk.clk
			audio_irq_irq             => irq_mapper_receiver0_irq,                                 --           audio_irq.irq
			audio_pll_ref_clk_clk     => audio_pll_ref_clk_clk,                                    --   audio_pll_ref_clk.clk
			audio_pll_ref_reset_reset => audio_pll_ref_reset_reset,                                -- audio_pll_ref_reset.reset
			audio_reset_reset         => open,                                                     --         audio_reset.reset
			audio_slave_address       => mm_interconnect_0_audio_subsystem_audio_slave_address,    --         audio_slave.address
			audio_slave_chipselect    => mm_interconnect_0_audio_subsystem_audio_slave_chipselect, --                    .chipselect
			audio_slave_read          => mm_interconnect_0_audio_subsystem_audio_slave_read,       --                    .read
			audio_slave_write         => mm_interconnect_0_audio_subsystem_audio_slave_write,      --                    .write
			audio_slave_writedata     => mm_interconnect_0_audio_subsystem_audio_slave_writedata,  --                    .writedata
			audio_slave_readdata      => mm_interconnect_0_audio_subsystem_audio_slave_readdata,   --                    .readdata
			sys_clk_clk               => system_pll_sys_clk_clk,                                   --             sys_clk.clk
			sys_reset_reset_n         => system_pll_reset_source_reset_ports_inv                   --           sys_reset.reset_n
		);

	camerad5m_0 : component nios_system_CameraD5M_0
		port map (
			camera_slave_readdata     => mm_interconnect_0_camerad5m_0_camera_slave_readdata, -- camera_slave.readdata
			clk_clk                   => system_pll_sys_clk_clk,                              --          clk.clk
			reset_reset_n             => system_pll_reset_source_reset_ports_inv,             --        reset.reset_n
			video_ext_PIXEL_CLK       => video_ext_1_PIXEL_CLK,                               --    video_ext.PIXEL_CLK
			video_ext_LINE_VALID      => video_ext_1_LINE_VALID,                              --             .LINE_VALID
			video_ext_FRAME_VALID     => video_ext_1_FRAME_VALID,                             --             .FRAME_VALID
			video_ext_pixel_clk_reset => video_ext_1_pixel_clk_reset,                         --             .pixel_clk_reset
			video_ext_PIXEL_DATA      => video_ext_1_PIXEL_DATA                               --             .PIXEL_DATA
		);

	expansion_jp5 : component nios_system_Expansion_JP5
		port map (
			clk        => system_pll_sys_clk_clk,                                                --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                        --                      reset.reset
			address    => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_readdata,   --                           .readdata
			GPIO       => expansion_jp5_export,                                                  --         external_interface.export
			irq        => irq_mapper_receiver1_irq                                               --                  interrupt.irq
		);

	flash : component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface
		generic map (
			FLASH_MEMORY_ADDRESS_WIDTH => 23
		)
		port map (
			i_avalon_chip_select       => mm_interconnect_0_flash_flash_data_chipselect,           --          flash_data.chipselect
			i_avalon_write             => mm_interconnect_0_flash_flash_data_write,                --                    .write
			i_avalon_read              => mm_interconnect_0_flash_flash_data_read,                 --                    .read
			i_avalon_address           => mm_interconnect_0_flash_flash_data_address,              --                    .address
			i_avalon_byteenable        => mm_interconnect_0_flash_flash_data_byteenable,           --                    .byteenable
			i_avalon_writedata         => mm_interconnect_0_flash_flash_data_writedata,            --                    .writedata
			o_avalon_readdata          => mm_interconnect_0_flash_flash_data_readdata,             --                    .readdata
			o_avalon_waitrequest       => mm_interconnect_0_flash_flash_data_waitrequest,          --                    .waitrequest
			i_clock                    => system_pll_sys_clk_clk,                                  --                 clk.clk
			i_reset_n                  => rst_controller_reset_out_reset_ports_inv,                --               reset.reset_n
			FL_ADDR                    => flash_ADDR,                                              --         conduit_end.export
			FL_CE_N                    => flash_CE_N,                                              --                    .export
			FL_OE_N                    => flash_OE_N,                                              --                    .export
			FL_WE_N                    => flash_WE_N,                                              --                    .export
			FL_RST_N                   => flash_RST_N,                                             --                    .export
			FL_DQ                      => flash_DQ,                                                --                    .export
			i_avalon_erase_write       => mm_interconnect_0_flash_flash_erase_control_write,       -- flash_erase_control.write
			i_avalon_erase_read        => mm_interconnect_0_flash_flash_erase_control_read,        --                    .read
			i_avalon_erase_byteenable  => mm_interconnect_0_flash_flash_erase_control_byteenable,  --                    .byteenable
			i_avalon_erase_writedata   => mm_interconnect_0_flash_flash_erase_control_writedata,   --                    .writedata
			i_avalon_erase_chip_select => mm_interconnect_0_flash_flash_erase_control_chipselect,  --                    .chipselect
			o_avalon_erase_readdata    => mm_interconnect_0_flash_flash_erase_control_readdata,    --                    .readdata
			o_avalon_erase_waitrequest => mm_interconnect_0_flash_flash_erase_control_waitrequest  --                    .waitrequest
		);

	green_leds : component nios_system_Green_LEDs
		port map (
			clk        => system_pll_sys_clk_clk,                                             --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                     --                      reset.reset
			address    => mm_interconnect_0_green_leds_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_green_leds_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_green_leds_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_green_leds_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_green_leds_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_green_leds_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_green_leds_avalon_parallel_port_slave_readdata,   --                           .readdata
			LEDG       => green_leds_export                                                   --         external_interface.export
		);

	interval_timer : component nios_system_Interval_Timer
		port map (
			clk        => system_pll_sys_clk_clk,                              --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => mm_interconnect_0_interval_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_interval_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_interval_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_interval_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_interval_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver4_irq                             --   irq.irq
		);

	jtag_uart : component nios_system_JTAG_UART
		port map (
			clk            => system_pll_sys_clk_clk,                                        --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver5_irq                                       --               irq.irq
		);

	jtag_uart_2nd_core : component nios_system_JTAG_UART
		port map (
			clk            => system_pll_sys_clk_clk,                                                 --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                               --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver5_irq                                            --               irq.irq
		);

	jtag_to_fpga_bridge : component nios_system_JTAG_to_FPGA_Bridge
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => system_pll_sys_clk_clk,                   --          clk.clk
			clk_reset_reset      => system_pll_reset_source_reset,            --    clk_reset.reset
			master_address       => jtag_to_fpga_bridge_master_address,       --       master.address
			master_readdata      => jtag_to_fpga_bridge_master_readdata,      --             .readdata
			master_read          => jtag_to_fpga_bridge_master_read,          --             .read
			master_write         => jtag_to_fpga_bridge_master_write,         --             .write
			master_writedata     => jtag_to_fpga_bridge_master_writedata,     --             .writedata
			master_waitrequest   => jtag_to_fpga_bridge_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_to_fpga_bridge_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_to_fpga_bridge_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                      -- master_reset.reset
		);

	nios2_floating_point : component fpoint_wrapper
		generic map (
			useDivider => 1
		)
		port map (
			clk    => processor1_custom_instruction_master_multi_slave_translator0_ci_master_clk,    -- s1.clk
			clk_en => processor1_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --   .clk_en
			dataa  => processor1_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  --   .dataa
			datab  => processor1_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --   .datab
			n      => processor1_custom_instruction_master_multi_slave_translator0_ci_master_n,      --   .n
			reset  => processor1_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --   .reset
			start  => processor1_custom_instruction_master_multi_slave_translator0_ci_master_start,  --   .start
			done   => processor1_custom_instruction_master_multi_slave_translator0_ci_master_done,   --   .done
			result => processor1_custom_instruction_master_multi_slave_translator0_ci_master_result  --   .result
		);

	nios2_floating_point_2nd_core : component fpoint_wrapper
		generic map (
			useDivider => 1
		)
		port map (
			clk    => processor2_custom_instruction_master_multi_slave_translator0_ci_master_clk,    -- s1.clk
			clk_en => processor2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --   .clk_en
			dataa  => processor2_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  --   .dataa
			datab  => processor2_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --   .datab
			n      => processor2_custom_instruction_master_multi_slave_translator0_ci_master_n,      --   .n
			reset  => processor2_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --   .reset
			start  => processor2_custom_instruction_master_multi_slave_translator0_ci_master_start,  --   .start
			done   => processor2_custom_instruction_master_multi_slave_translator0_ci_master_done,   --   .done
			result => processor2_custom_instruction_master_multi_slave_translator0_ci_master_result  --   .result
		);

	processor1 : component nios_system_Processor1
		port map (
			clk                                 => system_pll_sys_clk_clk,                                   --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                   --                          .reset_req
			d_address                           => processor1_data_master_address,                           --               data_master.address
			d_byteenable                        => processor1_data_master_byteenable,                        --                          .byteenable
			d_read                              => processor1_data_master_read,                              --                          .read
			d_readdata                          => processor1_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => processor1_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => processor1_data_master_write,                             --                          .write
			d_writedata                         => processor1_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => processor1_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => processor1_instruction_master_address,                    --        instruction_master.address
			i_read                              => processor1_instruction_master_read,                       --                          .read
			i_readdata                          => processor1_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => processor1_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => processor1_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => processor1_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_processor1_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_processor1_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_processor1_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_processor1_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_processor1_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_processor1_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_processor1_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_processor1_debug_mem_slave_writedata,   --                          .writedata
			E_ci_multi_done                     => processor1_custom_instruction_master_done,                -- custom_instruction_master.done
			E_ci_multi_clk_en                   => processor1_custom_instruction_master_clk_en,              --                          .clk_en
			E_ci_multi_start                    => processor1_custom_instruction_master_start,               --                          .start
			E_ci_result                         => processor1_custom_instruction_master_result,              --                          .result
			D_ci_a                              => processor1_custom_instruction_master_a,                   --                          .a
			D_ci_b                              => processor1_custom_instruction_master_b,                   --                          .b
			D_ci_c                              => processor1_custom_instruction_master_c,                   --                          .c
			D_ci_n                              => processor1_custom_instruction_master_n,                   --                          .n
			D_ci_readra                         => processor1_custom_instruction_master_readra,              --                          .readra
			D_ci_readrb                         => processor1_custom_instruction_master_readrb,              --                          .readrb
			D_ci_writerc                        => processor1_custom_instruction_master_writerc,             --                          .writerc
			E_ci_dataa                          => processor1_custom_instruction_master_dataa,               --                          .dataa
			E_ci_datab                          => processor1_custom_instruction_master_datab,               --                          .datab
			E_ci_multi_clock                    => processor1_custom_instruction_master_clk,                 --                          .clk
			E_ci_multi_reset                    => processor1_custom_instruction_master_reset,               --                          .reset
			E_ci_multi_reset_req                => processor1_custom_instruction_master_reset_req,           --                          .reset_req
			W_ci_estatus                        => processor1_custom_instruction_master_estatus,             --                          .estatus
			W_ci_ipending                       => processor1_custom_instruction_master_ipending             --                          .ipending
		);

	processor2 : component nios_system_Processor2
		port map (
			clk                                 => system_pll_sys_clk_clk,                                   --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,                   --                          .reset_req
			d_address                           => processor2_data_master_address,                           --               data_master.address
			d_byteenable                        => processor2_data_master_byteenable,                        --                          .byteenable
			d_read                              => processor2_data_master_read,                              --                          .read
			d_readdata                          => processor2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => processor2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => processor2_data_master_write,                             --                          .write
			d_writedata                         => processor2_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => processor2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => processor2_instruction_master_address,                    --        instruction_master.address
			i_read                              => processor2_instruction_master_read,                       --                          .read
			i_readdata                          => processor2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => processor2_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => processor2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => processor2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_processor2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_processor2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_processor2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_processor2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_processor2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_processor2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_processor2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_processor2_debug_mem_slave_writedata,   --                          .writedata
			E_ci_multi_done                     => processor2_custom_instruction_master_done,                -- custom_instruction_master.done
			E_ci_multi_clk_en                   => processor2_custom_instruction_master_clk_en,              --                          .clk_en
			E_ci_multi_start                    => processor2_custom_instruction_master_start,               --                          .start
			E_ci_result                         => processor2_custom_instruction_master_result,              --                          .result
			D_ci_a                              => processor2_custom_instruction_master_a,                   --                          .a
			D_ci_b                              => processor2_custom_instruction_master_b,                   --                          .b
			D_ci_c                              => processor2_custom_instruction_master_c,                   --                          .c
			D_ci_n                              => processor2_custom_instruction_master_n,                   --                          .n
			D_ci_readra                         => processor2_custom_instruction_master_readra,              --                          .readra
			D_ci_readrb                         => processor2_custom_instruction_master_readrb,              --                          .readrb
			D_ci_writerc                        => processor2_custom_instruction_master_writerc,             --                          .writerc
			E_ci_dataa                          => processor2_custom_instruction_master_dataa,               --                          .dataa
			E_ci_datab                          => processor2_custom_instruction_master_datab,               --                          .datab
			E_ci_multi_clock                    => processor2_custom_instruction_master_clk,                 --                          .clk
			E_ci_multi_reset                    => processor2_custom_instruction_master_reset,               --                          .reset
			E_ci_multi_reset_req                => processor2_custom_instruction_master_reset_req,           --                          .reset_req
			W_ci_estatus                        => processor2_custom_instruction_master_estatus,             --                          .estatus
			W_ci_ipending                       => processor2_custom_instruction_master_ipending             --                          .ipending
		);

	pushbuttons : component nios_system_Pushbuttons
		port map (
			clk        => system_pll_sys_clk_clk,                                              --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                      --                      reset.reset
			address    => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata,   --                           .readdata
			KEY        => pushbuttons_export,                                                  --         external_interface.export
			irq        => irq_mapper_receiver2_irq                                             --                  interrupt.irq
		);

	red_leds : component nios_system_Red_LEDs
		port map (
			clk        => system_pll_sys_clk_clk,                                           --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                   --                      reset.reset
			address    => mm_interconnect_0_red_leds_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_red_leds_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_red_leds_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_red_leds_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_red_leds_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_red_leds_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_red_leds_avalon_parallel_port_slave_readdata,   --                           .readdata
			LEDR       => red_leds_export                                                   --         external_interface.export
		);

	sdram : component nios_system_SDRAM
		port map (
			clk            => system_pll_sys_clk_clk,                          --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	sram : component nios_system_SRAM
		port map (
			clk           => system_pll_sys_clk_clk,                                 --                clk.clk
			reset         => rst_controller_reset_out_reset,                         --              reset.reset
			SRAM_DQ       => sram_DQ,                                                -- external_interface.export
			SRAM_ADDR     => sram_ADDR,                                              --                   .export
			SRAM_LB_N     => sram_LB_N,                                              --                   .export
			SRAM_UB_N     => sram_UB_N,                                              --                   .export
			SRAM_CE_N     => sram_CE_N,                                              --                   .export
			SRAM_OE_N     => sram_OE_N,                                              --                   .export
			SRAM_WE_N     => sram_WE_N,                                              --                   .export
			address       => mm_interconnect_0_sram_avalon_sram_slave_address,       --  avalon_sram_slave.address
			byteenable    => mm_interconnect_0_sram_avalon_sram_slave_byteenable,    --                   .byteenable
			read          => mm_interconnect_0_sram_avalon_sram_slave_read,          --                   .read
			write         => mm_interconnect_0_sram_avalon_sram_slave_write,         --                   .write
			writedata     => mm_interconnect_0_sram_avalon_sram_slave_writedata,     --                   .writedata
			readdata      => mm_interconnect_0_sram_avalon_sram_slave_readdata,      --                   .readdata
			readdatavalid => mm_interconnect_0_sram_avalon_sram_slave_readdatavalid  --                   .readdatavalid
		);

	serial_port : component nios_system_Serial_Port
		port map (
			clk        => system_pll_sys_clk_clk,                                      --                clk.clk
			reset      => rst_controller_reset_out_reset,                              --              reset.reset
			address    => mm_interconnect_0_serial_port_avalon_rs232_slave_address(0), -- avalon_rs232_slave.address
			chipselect => mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect, --                   .chipselect
			byteenable => mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable, --                   .byteenable
			read       => mm_interconnect_0_serial_port_avalon_rs232_slave_read,       --                   .read
			write      => mm_interconnect_0_serial_port_avalon_rs232_slave_write,      --                   .write
			writedata  => mm_interconnect_0_serial_port_avalon_rs232_slave_writedata,  --                   .writedata
			readdata   => mm_interconnect_0_serial_port_avalon_rs232_slave_readdata,   --                   .readdata
			irq        => irq_mapper_receiver3_irq,                                    --          interrupt.irq
			UART_RXD   => serial_port_RXD,                                             -- external_interface.export
			UART_TXD   => serial_port_TXD                                              --                   .export
		);

	slider_switches : component nios_system_Slider_Switches
		port map (
			clk        => system_pll_sys_clk_clk,                                                  --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                          --                      reset.reset
			address    => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_readdata,   --                           .readdata
			SW         => slider_switches_export                                                   --         external_interface.export
		);

	sysid : component nios_system_SysID
		port map (
			clock    => system_pll_sys_clk_clk,                           --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	system_pll : component nios_system_System_PLL
		port map (
			ref_clk_clk        => system_pll_ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => system_pll_ref_reset_reset,    --    ref_reset.reset
			sys_clk_clk        => system_pll_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                 --    sdram_clk.clk
			reset_source_reset => system_pll_reset_source_reset  -- reset_source.reset
		);

	processor1_custom_instruction_master_translator : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 1
		)
		port map (
			ci_slave_dataa            => processor1_custom_instruction_master_dataa,                                --        ci_slave.dataa
			ci_slave_datab            => processor1_custom_instruction_master_datab,                                --                .datab
			ci_slave_result           => processor1_custom_instruction_master_result,                               --                .result
			ci_slave_n                => processor1_custom_instruction_master_n,                                    --                .n
			ci_slave_readra           => processor1_custom_instruction_master_readra,                               --                .readra
			ci_slave_readrb           => processor1_custom_instruction_master_readrb,                               --                .readrb
			ci_slave_writerc          => processor1_custom_instruction_master_writerc,                              --                .writerc
			ci_slave_a                => processor1_custom_instruction_master_a,                                    --                .a
			ci_slave_b                => processor1_custom_instruction_master_b,                                    --                .b
			ci_slave_c                => processor1_custom_instruction_master_c,                                    --                .c
			ci_slave_ipending         => processor1_custom_instruction_master_ipending,                             --                .ipending
			ci_slave_estatus          => processor1_custom_instruction_master_estatus,                              --                .estatus
			ci_slave_multi_clk        => processor1_custom_instruction_master_clk,                                  --                .clk
			ci_slave_multi_reset      => processor1_custom_instruction_master_reset,                                --                .reset
			ci_slave_multi_clken      => processor1_custom_instruction_master_clk_en,                               --                .clk_en
			ci_slave_multi_reset_req  => processor1_custom_instruction_master_reset_req,                            --                .reset_req
			ci_slave_multi_start      => processor1_custom_instruction_master_start,                                --                .start
			ci_slave_multi_done       => processor1_custom_instruction_master_done,                                 --                .done
			comb_ci_master_dataa      => open,                                                                      --  comb_ci_master.dataa
			comb_ci_master_datab      => open,                                                                      --                .datab
			comb_ci_master_result     => open,                                                                      --                .result
			comb_ci_master_n          => open,                                                                      --                .n
			comb_ci_master_readra     => open,                                                                      --                .readra
			comb_ci_master_readrb     => open,                                                                      --                .readrb
			comb_ci_master_writerc    => open,                                                                      --                .writerc
			comb_ci_master_a          => open,                                                                      --                .a
			comb_ci_master_b          => open,                                                                      --                .b
			comb_ci_master_c          => open,                                                                      --                .c
			comb_ci_master_ipending   => open,                                                                      --                .ipending
			comb_ci_master_estatus    => open,                                                                      --                .estatus
			multi_ci_master_clk       => processor1_custom_instruction_master_translator_multi_ci_master_clk,       -- multi_ci_master.clk
			multi_ci_master_reset     => processor1_custom_instruction_master_translator_multi_ci_master_reset,     --                .reset
			multi_ci_master_clken     => processor1_custom_instruction_master_translator_multi_ci_master_clk_en,    --                .clk_en
			multi_ci_master_reset_req => processor1_custom_instruction_master_translator_multi_ci_master_reset_req, --                .reset_req
			multi_ci_master_start     => processor1_custom_instruction_master_translator_multi_ci_master_start,     --                .start
			multi_ci_master_done      => processor1_custom_instruction_master_translator_multi_ci_master_done,      --                .done
			multi_ci_master_dataa     => processor1_custom_instruction_master_translator_multi_ci_master_dataa,     --                .dataa
			multi_ci_master_datab     => processor1_custom_instruction_master_translator_multi_ci_master_datab,     --                .datab
			multi_ci_master_result    => processor1_custom_instruction_master_translator_multi_ci_master_result,    --                .result
			multi_ci_master_n         => processor1_custom_instruction_master_translator_multi_ci_master_n,         --                .n
			multi_ci_master_readra    => processor1_custom_instruction_master_translator_multi_ci_master_readra,    --                .readra
			multi_ci_master_readrb    => processor1_custom_instruction_master_translator_multi_ci_master_readrb,    --                .readrb
			multi_ci_master_writerc   => processor1_custom_instruction_master_translator_multi_ci_master_writerc,   --                .writerc
			multi_ci_master_a         => processor1_custom_instruction_master_translator_multi_ci_master_a,         --                .a
			multi_ci_master_b         => processor1_custom_instruction_master_translator_multi_ci_master_b,         --                .b
			multi_ci_master_c         => processor1_custom_instruction_master_translator_multi_ci_master_c,         --                .c
			ci_slave_multi_dataa      => "00000000000000000000000000000000",                                        --     (terminated)
			ci_slave_multi_datab      => "00000000000000000000000000000000",                                        --     (terminated)
			ci_slave_multi_result     => open,                                                                      --     (terminated)
			ci_slave_multi_n          => "00000000",                                                                --     (terminated)
			ci_slave_multi_readra     => '0',                                                                       --     (terminated)
			ci_slave_multi_readrb     => '0',                                                                       --     (terminated)
			ci_slave_multi_writerc    => '0',                                                                       --     (terminated)
			ci_slave_multi_a          => "00000",                                                                   --     (terminated)
			ci_slave_multi_b          => "00000",                                                                   --     (terminated)
			ci_slave_multi_c          => "00000"                                                                    --     (terminated)
		);

	processor1_custom_instruction_master_multi_xconnect : component nios_system_Processor1_custom_instruction_master_multi_xconnect
		port map (
			ci_slave_dataa       => processor1_custom_instruction_master_translator_multi_ci_master_dataa,     --   ci_slave.dataa
			ci_slave_datab       => processor1_custom_instruction_master_translator_multi_ci_master_datab,     --           .datab
			ci_slave_result      => processor1_custom_instruction_master_translator_multi_ci_master_result,    --           .result
			ci_slave_n           => processor1_custom_instruction_master_translator_multi_ci_master_n,         --           .n
			ci_slave_readra      => processor1_custom_instruction_master_translator_multi_ci_master_readra,    --           .readra
			ci_slave_readrb      => processor1_custom_instruction_master_translator_multi_ci_master_readrb,    --           .readrb
			ci_slave_writerc     => processor1_custom_instruction_master_translator_multi_ci_master_writerc,   --           .writerc
			ci_slave_a           => processor1_custom_instruction_master_translator_multi_ci_master_a,         --           .a
			ci_slave_b           => processor1_custom_instruction_master_translator_multi_ci_master_b,         --           .b
			ci_slave_c           => processor1_custom_instruction_master_translator_multi_ci_master_c,         --           .c
			ci_slave_ipending    => open,                                                                      --           .ipending
			ci_slave_estatus     => open,                                                                      --           .estatus
			ci_slave_clk         => processor1_custom_instruction_master_translator_multi_ci_master_clk,       --           .clk
			ci_slave_reset       => processor1_custom_instruction_master_translator_multi_ci_master_reset,     --           .reset
			ci_slave_clken       => processor1_custom_instruction_master_translator_multi_ci_master_clk_en,    --           .clk_en
			ci_slave_reset_req   => processor1_custom_instruction_master_translator_multi_ci_master_reset_req, --           .reset_req
			ci_slave_start       => processor1_custom_instruction_master_translator_multi_ci_master_start,     --           .start
			ci_slave_done        => processor1_custom_instruction_master_translator_multi_ci_master_done,      --           .done
			ci_master0_dataa     => processor1_custom_instruction_master_multi_xconnect_ci_master0_dataa,      -- ci_master0.dataa
			ci_master0_datab     => processor1_custom_instruction_master_multi_xconnect_ci_master0_datab,      --           .datab
			ci_master0_result    => processor1_custom_instruction_master_multi_xconnect_ci_master0_result,     --           .result
			ci_master0_n         => processor1_custom_instruction_master_multi_xconnect_ci_master0_n,          --           .n
			ci_master0_readra    => processor1_custom_instruction_master_multi_xconnect_ci_master0_readra,     --           .readra
			ci_master0_readrb    => processor1_custom_instruction_master_multi_xconnect_ci_master0_readrb,     --           .readrb
			ci_master0_writerc   => processor1_custom_instruction_master_multi_xconnect_ci_master0_writerc,    --           .writerc
			ci_master0_a         => processor1_custom_instruction_master_multi_xconnect_ci_master0_a,          --           .a
			ci_master0_b         => processor1_custom_instruction_master_multi_xconnect_ci_master0_b,          --           .b
			ci_master0_c         => processor1_custom_instruction_master_multi_xconnect_ci_master0_c,          --           .c
			ci_master0_ipending  => processor1_custom_instruction_master_multi_xconnect_ci_master0_ipending,   --           .ipending
			ci_master0_estatus   => processor1_custom_instruction_master_multi_xconnect_ci_master0_estatus,    --           .estatus
			ci_master0_clk       => processor1_custom_instruction_master_multi_xconnect_ci_master0_clk,        --           .clk
			ci_master0_reset     => processor1_custom_instruction_master_multi_xconnect_ci_master0_reset,      --           .reset
			ci_master0_clken     => processor1_custom_instruction_master_multi_xconnect_ci_master0_clk_en,     --           .clk_en
			ci_master0_reset_req => processor1_custom_instruction_master_multi_xconnect_ci_master0_reset_req,  --           .reset_req
			ci_master0_start     => processor1_custom_instruction_master_multi_xconnect_ci_master0_start,      --           .start
			ci_master0_done      => processor1_custom_instruction_master_multi_xconnect_ci_master0_done        --           .done
		);

	processor1_custom_instruction_master_multi_slave_translator0 : component altera_customins_slave_translator
		generic map (
			N_WIDTH          => 2,
			USE_DONE         => 1,
			NUM_FIXED_CYCLES => 1
		)
		port map (
			ci_slave_dataa      => processor1_custom_instruction_master_multi_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab      => processor1_custom_instruction_master_multi_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result     => processor1_custom_instruction_master_multi_xconnect_ci_master0_result,         --          .result
			ci_slave_n          => processor1_custom_instruction_master_multi_xconnect_ci_master0_n,              --          .n
			ci_slave_readra     => processor1_custom_instruction_master_multi_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb     => processor1_custom_instruction_master_multi_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc    => processor1_custom_instruction_master_multi_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a          => processor1_custom_instruction_master_multi_xconnect_ci_master0_a,              --          .a
			ci_slave_b          => processor1_custom_instruction_master_multi_xconnect_ci_master0_b,              --          .b
			ci_slave_c          => processor1_custom_instruction_master_multi_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending   => processor1_custom_instruction_master_multi_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus    => processor1_custom_instruction_master_multi_xconnect_ci_master0_estatus,        --          .estatus
			ci_slave_clk        => processor1_custom_instruction_master_multi_xconnect_ci_master0_clk,            --          .clk
			ci_slave_clken      => processor1_custom_instruction_master_multi_xconnect_ci_master0_clk_en,         --          .clk_en
			ci_slave_reset_req  => processor1_custom_instruction_master_multi_xconnect_ci_master0_reset_req,      --          .reset_req
			ci_slave_reset      => processor1_custom_instruction_master_multi_xconnect_ci_master0_reset,          --          .reset
			ci_slave_start      => processor1_custom_instruction_master_multi_xconnect_ci_master0_start,          --          .start
			ci_slave_done       => processor1_custom_instruction_master_multi_xconnect_ci_master0_done,           --          .done
			ci_master_dataa     => processor1_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab     => processor1_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --          .datab
			ci_master_result    => processor1_custom_instruction_master_multi_slave_translator0_ci_master_result, --          .result
			ci_master_n         => processor1_custom_instruction_master_multi_slave_translator0_ci_master_n,      --          .n
			ci_master_clk       => processor1_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --          .clk
			ci_master_clken     => processor1_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --          .clk_en
			ci_master_reset     => processor1_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --          .reset
			ci_master_start     => processor1_custom_instruction_master_multi_slave_translator0_ci_master_start,  --          .start
			ci_master_done      => processor1_custom_instruction_master_multi_slave_translator0_ci_master_done,   --          .done
			ci_master_readra    => open,                                                                          -- (terminated)
			ci_master_readrb    => open,                                                                          -- (terminated)
			ci_master_writerc   => open,                                                                          -- (terminated)
			ci_master_a         => open,                                                                          -- (terminated)
			ci_master_b         => open,                                                                          -- (terminated)
			ci_master_c         => open,                                                                          -- (terminated)
			ci_master_ipending  => open,                                                                          -- (terminated)
			ci_master_estatus   => open,                                                                          -- (terminated)
			ci_master_reset_req => open                                                                           -- (terminated)
		);

	processor2_custom_instruction_master_translator : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 1
		)
		port map (
			ci_slave_dataa            => processor2_custom_instruction_master_dataa,                                --        ci_slave.dataa
			ci_slave_datab            => processor2_custom_instruction_master_datab,                                --                .datab
			ci_slave_result           => processor2_custom_instruction_master_result,                               --                .result
			ci_slave_n                => processor2_custom_instruction_master_n,                                    --                .n
			ci_slave_readra           => processor2_custom_instruction_master_readra,                               --                .readra
			ci_slave_readrb           => processor2_custom_instruction_master_readrb,                               --                .readrb
			ci_slave_writerc          => processor2_custom_instruction_master_writerc,                              --                .writerc
			ci_slave_a                => processor2_custom_instruction_master_a,                                    --                .a
			ci_slave_b                => processor2_custom_instruction_master_b,                                    --                .b
			ci_slave_c                => processor2_custom_instruction_master_c,                                    --                .c
			ci_slave_ipending         => processor2_custom_instruction_master_ipending,                             --                .ipending
			ci_slave_estatus          => processor2_custom_instruction_master_estatus,                              --                .estatus
			ci_slave_multi_clk        => processor2_custom_instruction_master_clk,                                  --                .clk
			ci_slave_multi_reset      => processor2_custom_instruction_master_reset,                                --                .reset
			ci_slave_multi_clken      => processor2_custom_instruction_master_clk_en,                               --                .clk_en
			ci_slave_multi_reset_req  => processor2_custom_instruction_master_reset_req,                            --                .reset_req
			ci_slave_multi_start      => processor2_custom_instruction_master_start,                                --                .start
			ci_slave_multi_done       => processor2_custom_instruction_master_done,                                 --                .done
			comb_ci_master_dataa      => open,                                                                      --  comb_ci_master.dataa
			comb_ci_master_datab      => open,                                                                      --                .datab
			comb_ci_master_result     => open,                                                                      --                .result
			comb_ci_master_n          => open,                                                                      --                .n
			comb_ci_master_readra     => open,                                                                      --                .readra
			comb_ci_master_readrb     => open,                                                                      --                .readrb
			comb_ci_master_writerc    => open,                                                                      --                .writerc
			comb_ci_master_a          => open,                                                                      --                .a
			comb_ci_master_b          => open,                                                                      --                .b
			comb_ci_master_c          => open,                                                                      --                .c
			comb_ci_master_ipending   => open,                                                                      --                .ipending
			comb_ci_master_estatus    => open,                                                                      --                .estatus
			multi_ci_master_clk       => processor2_custom_instruction_master_translator_multi_ci_master_clk,       -- multi_ci_master.clk
			multi_ci_master_reset     => processor2_custom_instruction_master_translator_multi_ci_master_reset,     --                .reset
			multi_ci_master_clken     => processor2_custom_instruction_master_translator_multi_ci_master_clk_en,    --                .clk_en
			multi_ci_master_reset_req => processor2_custom_instruction_master_translator_multi_ci_master_reset_req, --                .reset_req
			multi_ci_master_start     => processor2_custom_instruction_master_translator_multi_ci_master_start,     --                .start
			multi_ci_master_done      => processor2_custom_instruction_master_translator_multi_ci_master_done,      --                .done
			multi_ci_master_dataa     => processor2_custom_instruction_master_translator_multi_ci_master_dataa,     --                .dataa
			multi_ci_master_datab     => processor2_custom_instruction_master_translator_multi_ci_master_datab,     --                .datab
			multi_ci_master_result    => processor2_custom_instruction_master_translator_multi_ci_master_result,    --                .result
			multi_ci_master_n         => processor2_custom_instruction_master_translator_multi_ci_master_n,         --                .n
			multi_ci_master_readra    => processor2_custom_instruction_master_translator_multi_ci_master_readra,    --                .readra
			multi_ci_master_readrb    => processor2_custom_instruction_master_translator_multi_ci_master_readrb,    --                .readrb
			multi_ci_master_writerc   => processor2_custom_instruction_master_translator_multi_ci_master_writerc,   --                .writerc
			multi_ci_master_a         => processor2_custom_instruction_master_translator_multi_ci_master_a,         --                .a
			multi_ci_master_b         => processor2_custom_instruction_master_translator_multi_ci_master_b,         --                .b
			multi_ci_master_c         => processor2_custom_instruction_master_translator_multi_ci_master_c,         --                .c
			ci_slave_multi_dataa      => "00000000000000000000000000000000",                                        --     (terminated)
			ci_slave_multi_datab      => "00000000000000000000000000000000",                                        --     (terminated)
			ci_slave_multi_result     => open,                                                                      --     (terminated)
			ci_slave_multi_n          => "00000000",                                                                --     (terminated)
			ci_slave_multi_readra     => '0',                                                                       --     (terminated)
			ci_slave_multi_readrb     => '0',                                                                       --     (terminated)
			ci_slave_multi_writerc    => '0',                                                                       --     (terminated)
			ci_slave_multi_a          => "00000",                                                                   --     (terminated)
			ci_slave_multi_b          => "00000",                                                                   --     (terminated)
			ci_slave_multi_c          => "00000"                                                                    --     (terminated)
		);

	processor2_custom_instruction_master_multi_xconnect : component nios_system_Processor1_custom_instruction_master_multi_xconnect
		port map (
			ci_slave_dataa       => processor2_custom_instruction_master_translator_multi_ci_master_dataa,     --   ci_slave.dataa
			ci_slave_datab       => processor2_custom_instruction_master_translator_multi_ci_master_datab,     --           .datab
			ci_slave_result      => processor2_custom_instruction_master_translator_multi_ci_master_result,    --           .result
			ci_slave_n           => processor2_custom_instruction_master_translator_multi_ci_master_n,         --           .n
			ci_slave_readra      => processor2_custom_instruction_master_translator_multi_ci_master_readra,    --           .readra
			ci_slave_readrb      => processor2_custom_instruction_master_translator_multi_ci_master_readrb,    --           .readrb
			ci_slave_writerc     => processor2_custom_instruction_master_translator_multi_ci_master_writerc,   --           .writerc
			ci_slave_a           => processor2_custom_instruction_master_translator_multi_ci_master_a,         --           .a
			ci_slave_b           => processor2_custom_instruction_master_translator_multi_ci_master_b,         --           .b
			ci_slave_c           => processor2_custom_instruction_master_translator_multi_ci_master_c,         --           .c
			ci_slave_ipending    => open,                                                                      --           .ipending
			ci_slave_estatus     => open,                                                                      --           .estatus
			ci_slave_clk         => processor2_custom_instruction_master_translator_multi_ci_master_clk,       --           .clk
			ci_slave_reset       => processor2_custom_instruction_master_translator_multi_ci_master_reset,     --           .reset
			ci_slave_clken       => processor2_custom_instruction_master_translator_multi_ci_master_clk_en,    --           .clk_en
			ci_slave_reset_req   => processor2_custom_instruction_master_translator_multi_ci_master_reset_req, --           .reset_req
			ci_slave_start       => processor2_custom_instruction_master_translator_multi_ci_master_start,     --           .start
			ci_slave_done        => processor2_custom_instruction_master_translator_multi_ci_master_done,      --           .done
			ci_master0_dataa     => processor2_custom_instruction_master_multi_xconnect_ci_master0_dataa,      -- ci_master0.dataa
			ci_master0_datab     => processor2_custom_instruction_master_multi_xconnect_ci_master0_datab,      --           .datab
			ci_master0_result    => processor2_custom_instruction_master_multi_xconnect_ci_master0_result,     --           .result
			ci_master0_n         => processor2_custom_instruction_master_multi_xconnect_ci_master0_n,          --           .n
			ci_master0_readra    => processor2_custom_instruction_master_multi_xconnect_ci_master0_readra,     --           .readra
			ci_master0_readrb    => processor2_custom_instruction_master_multi_xconnect_ci_master0_readrb,     --           .readrb
			ci_master0_writerc   => processor2_custom_instruction_master_multi_xconnect_ci_master0_writerc,    --           .writerc
			ci_master0_a         => processor2_custom_instruction_master_multi_xconnect_ci_master0_a,          --           .a
			ci_master0_b         => processor2_custom_instruction_master_multi_xconnect_ci_master0_b,          --           .b
			ci_master0_c         => processor2_custom_instruction_master_multi_xconnect_ci_master0_c,          --           .c
			ci_master0_ipending  => processor2_custom_instruction_master_multi_xconnect_ci_master0_ipending,   --           .ipending
			ci_master0_estatus   => processor2_custom_instruction_master_multi_xconnect_ci_master0_estatus,    --           .estatus
			ci_master0_clk       => processor2_custom_instruction_master_multi_xconnect_ci_master0_clk,        --           .clk
			ci_master0_reset     => processor2_custom_instruction_master_multi_xconnect_ci_master0_reset,      --           .reset
			ci_master0_clken     => processor2_custom_instruction_master_multi_xconnect_ci_master0_clk_en,     --           .clk_en
			ci_master0_reset_req => processor2_custom_instruction_master_multi_xconnect_ci_master0_reset_req,  --           .reset_req
			ci_master0_start     => processor2_custom_instruction_master_multi_xconnect_ci_master0_start,      --           .start
			ci_master0_done      => processor2_custom_instruction_master_multi_xconnect_ci_master0_done        --           .done
		);

	processor2_custom_instruction_master_multi_slave_translator0 : component altera_customins_slave_translator
		generic map (
			N_WIDTH          => 2,
			USE_DONE         => 1,
			NUM_FIXED_CYCLES => 1
		)
		port map (
			ci_slave_dataa      => processor2_custom_instruction_master_multi_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab      => processor2_custom_instruction_master_multi_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result     => processor2_custom_instruction_master_multi_xconnect_ci_master0_result,         --          .result
			ci_slave_n          => processor2_custom_instruction_master_multi_xconnect_ci_master0_n,              --          .n
			ci_slave_readra     => processor2_custom_instruction_master_multi_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb     => processor2_custom_instruction_master_multi_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc    => processor2_custom_instruction_master_multi_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a          => processor2_custom_instruction_master_multi_xconnect_ci_master0_a,              --          .a
			ci_slave_b          => processor2_custom_instruction_master_multi_xconnect_ci_master0_b,              --          .b
			ci_slave_c          => processor2_custom_instruction_master_multi_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending   => processor2_custom_instruction_master_multi_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus    => processor2_custom_instruction_master_multi_xconnect_ci_master0_estatus,        --          .estatus
			ci_slave_clk        => processor2_custom_instruction_master_multi_xconnect_ci_master0_clk,            --          .clk
			ci_slave_clken      => processor2_custom_instruction_master_multi_xconnect_ci_master0_clk_en,         --          .clk_en
			ci_slave_reset_req  => processor2_custom_instruction_master_multi_xconnect_ci_master0_reset_req,      --          .reset_req
			ci_slave_reset      => processor2_custom_instruction_master_multi_xconnect_ci_master0_reset,          --          .reset
			ci_slave_start      => processor2_custom_instruction_master_multi_xconnect_ci_master0_start,          --          .start
			ci_slave_done       => processor2_custom_instruction_master_multi_xconnect_ci_master0_done,           --          .done
			ci_master_dataa     => processor2_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab     => processor2_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --          .datab
			ci_master_result    => processor2_custom_instruction_master_multi_slave_translator0_ci_master_result, --          .result
			ci_master_n         => processor2_custom_instruction_master_multi_slave_translator0_ci_master_n,      --          .n
			ci_master_clk       => processor2_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --          .clk
			ci_master_clken     => processor2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --          .clk_en
			ci_master_reset     => processor2_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --          .reset
			ci_master_start     => processor2_custom_instruction_master_multi_slave_translator0_ci_master_start,  --          .start
			ci_master_done      => processor2_custom_instruction_master_multi_slave_translator0_ci_master_done,   --          .done
			ci_master_readra    => open,                                                                          -- (terminated)
			ci_master_readrb    => open,                                                                          -- (terminated)
			ci_master_writerc   => open,                                                                          -- (terminated)
			ci_master_a         => open,                                                                          -- (terminated)
			ci_master_b         => open,                                                                          -- (terminated)
			ci_master_c         => open,                                                                          -- (terminated)
			ci_master_ipending  => open,                                                                          -- (terminated)
			ci_master_estatus   => open,                                                                          -- (terminated)
			ci_master_reset_req => open                                                                           -- (terminated)
		);

	mm_interconnect_0 : component nios_system_mm_interconnect_0
		port map (
			System_PLL_sys_clk_clk                                    => system_pll_sys_clk_clk,                                                  --                                  System_PLL_sys_clk.clk
			JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                          -- JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset.reset
			JTAG_UART_2nd_Core_reset_reset_bridge_in_reset_reset      => rst_controller_reset_out_reset,                                          --      JTAG_UART_2nd_Core_reset_reset_bridge_in_reset.reset
			Processor1_reset_reset_bridge_in_reset_reset              => rst_controller_001_reset_out_reset,                                      --              Processor1_reset_reset_bridge_in_reset.reset
			Processor2_reset_reset_bridge_in_reset_reset              => rst_controller_002_reset_out_reset,                                      --              Processor2_reset_reset_bridge_in_reset.reset
			JTAG_to_FPGA_Bridge_master_address                        => jtag_to_fpga_bridge_master_address,                                      --                          JTAG_to_FPGA_Bridge_master.address
			JTAG_to_FPGA_Bridge_master_waitrequest                    => jtag_to_fpga_bridge_master_waitrequest,                                  --                                                    .waitrequest
			JTAG_to_FPGA_Bridge_master_byteenable                     => jtag_to_fpga_bridge_master_byteenable,                                   --                                                    .byteenable
			JTAG_to_FPGA_Bridge_master_read                           => jtag_to_fpga_bridge_master_read,                                         --                                                    .read
			JTAG_to_FPGA_Bridge_master_readdata                       => jtag_to_fpga_bridge_master_readdata,                                     --                                                    .readdata
			JTAG_to_FPGA_Bridge_master_readdatavalid                  => jtag_to_fpga_bridge_master_readdatavalid,                                --                                                    .readdatavalid
			JTAG_to_FPGA_Bridge_master_write                          => jtag_to_fpga_bridge_master_write,                                        --                                                    .write
			JTAG_to_FPGA_Bridge_master_writedata                      => jtag_to_fpga_bridge_master_writedata,                                    --                                                    .writedata
			Processor1_data_master_address                            => processor1_data_master_address,                                          --                              Processor1_data_master.address
			Processor1_data_master_waitrequest                        => processor1_data_master_waitrequest,                                      --                                                    .waitrequest
			Processor1_data_master_byteenable                         => processor1_data_master_byteenable,                                       --                                                    .byteenable
			Processor1_data_master_read                               => processor1_data_master_read,                                             --                                                    .read
			Processor1_data_master_readdata                           => processor1_data_master_readdata,                                         --                                                    .readdata
			Processor1_data_master_write                              => processor1_data_master_write,                                            --                                                    .write
			Processor1_data_master_writedata                          => processor1_data_master_writedata,                                        --                                                    .writedata
			Processor1_data_master_debugaccess                        => processor1_data_master_debugaccess,                                      --                                                    .debugaccess
			Processor1_instruction_master_address                     => processor1_instruction_master_address,                                   --                       Processor1_instruction_master.address
			Processor1_instruction_master_waitrequest                 => processor1_instruction_master_waitrequest,                               --                                                    .waitrequest
			Processor1_instruction_master_read                        => processor1_instruction_master_read,                                      --                                                    .read
			Processor1_instruction_master_readdata                    => processor1_instruction_master_readdata,                                  --                                                    .readdata
			Processor2_data_master_address                            => processor2_data_master_address,                                          --                              Processor2_data_master.address
			Processor2_data_master_waitrequest                        => processor2_data_master_waitrequest,                                      --                                                    .waitrequest
			Processor2_data_master_byteenable                         => processor2_data_master_byteenable,                                       --                                                    .byteenable
			Processor2_data_master_read                               => processor2_data_master_read,                                             --                                                    .read
			Processor2_data_master_readdata                           => processor2_data_master_readdata,                                         --                                                    .readdata
			Processor2_data_master_write                              => processor2_data_master_write,                                            --                                                    .write
			Processor2_data_master_writedata                          => processor2_data_master_writedata,                                        --                                                    .writedata
			Processor2_data_master_debugaccess                        => processor2_data_master_debugaccess,                                      --                                                    .debugaccess
			Processor2_instruction_master_address                     => processor2_instruction_master_address,                                   --                       Processor2_instruction_master.address
			Processor2_instruction_master_waitrequest                 => processor2_instruction_master_waitrequest,                               --                                                    .waitrequest
			Processor2_instruction_master_read                        => processor2_instruction_master_read,                                      --                                                    .read
			Processor2_instruction_master_readdata                    => processor2_instruction_master_readdata,                                  --                                                    .readdata
			Audio_Subsystem_audio_slave_address                       => mm_interconnect_0_audio_subsystem_audio_slave_address,                   --                         Audio_Subsystem_audio_slave.address
			Audio_Subsystem_audio_slave_write                         => mm_interconnect_0_audio_subsystem_audio_slave_write,                     --                                                    .write
			Audio_Subsystem_audio_slave_read                          => mm_interconnect_0_audio_subsystem_audio_slave_read,                      --                                                    .read
			Audio_Subsystem_audio_slave_readdata                      => mm_interconnect_0_audio_subsystem_audio_slave_readdata,                  --                                                    .readdata
			Audio_Subsystem_audio_slave_writedata                     => mm_interconnect_0_audio_subsystem_audio_slave_writedata,                 --                                                    .writedata
			Audio_Subsystem_audio_slave_chipselect                    => mm_interconnect_0_audio_subsystem_audio_slave_chipselect,                --                                                    .chipselect
			AV_Config_avalon_av_config_slave_address                  => mm_interconnect_0_av_config_avalon_av_config_slave_address,              --                    AV_Config_avalon_av_config_slave.address
			AV_Config_avalon_av_config_slave_write                    => mm_interconnect_0_av_config_avalon_av_config_slave_write,                --                                                    .write
			AV_Config_avalon_av_config_slave_read                     => mm_interconnect_0_av_config_avalon_av_config_slave_read,                 --                                                    .read
			AV_Config_avalon_av_config_slave_readdata                 => mm_interconnect_0_av_config_avalon_av_config_slave_readdata,             --                                                    .readdata
			AV_Config_avalon_av_config_slave_writedata                => mm_interconnect_0_av_config_avalon_av_config_slave_writedata,            --                                                    .writedata
			AV_Config_avalon_av_config_slave_byteenable               => mm_interconnect_0_av_config_avalon_av_config_slave_byteenable,           --                                                    .byteenable
			AV_Config_avalon_av_config_slave_waitrequest              => mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest,          --                                                    .waitrequest
			CameraD5M_0_camera_slave_readdata                         => mm_interconnect_0_camerad5m_0_camera_slave_readdata,                     --                            CameraD5M_0_camera_slave.readdata
			Expansion_JP5_avalon_parallel_port_slave_address          => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_address,      --            Expansion_JP5_avalon_parallel_port_slave.address
			Expansion_JP5_avalon_parallel_port_slave_write            => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_write,        --                                                    .write
			Expansion_JP5_avalon_parallel_port_slave_read             => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_read,         --                                                    .read
			Expansion_JP5_avalon_parallel_port_slave_readdata         => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_readdata,     --                                                    .readdata
			Expansion_JP5_avalon_parallel_port_slave_writedata        => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_writedata,    --                                                    .writedata
			Expansion_JP5_avalon_parallel_port_slave_byteenable       => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_byteenable,   --                                                    .byteenable
			Expansion_JP5_avalon_parallel_port_slave_chipselect       => mm_interconnect_0_expansion_jp5_avalon_parallel_port_slave_chipselect,   --                                                    .chipselect
			Flash_flash_data_address                                  => mm_interconnect_0_flash_flash_data_address,                              --                                    Flash_flash_data.address
			Flash_flash_data_write                                    => mm_interconnect_0_flash_flash_data_write,                                --                                                    .write
			Flash_flash_data_read                                     => mm_interconnect_0_flash_flash_data_read,                                 --                                                    .read
			Flash_flash_data_readdata                                 => mm_interconnect_0_flash_flash_data_readdata,                             --                                                    .readdata
			Flash_flash_data_writedata                                => mm_interconnect_0_flash_flash_data_writedata,                            --                                                    .writedata
			Flash_flash_data_byteenable                               => mm_interconnect_0_flash_flash_data_byteenable,                           --                                                    .byteenable
			Flash_flash_data_waitrequest                              => mm_interconnect_0_flash_flash_data_waitrequest,                          --                                                    .waitrequest
			Flash_flash_data_chipselect                               => mm_interconnect_0_flash_flash_data_chipselect,                           --                                                    .chipselect
			Flash_flash_erase_control_write                           => mm_interconnect_0_flash_flash_erase_control_write,                       --                           Flash_flash_erase_control.write
			Flash_flash_erase_control_read                            => mm_interconnect_0_flash_flash_erase_control_read,                        --                                                    .read
			Flash_flash_erase_control_readdata                        => mm_interconnect_0_flash_flash_erase_control_readdata,                    --                                                    .readdata
			Flash_flash_erase_control_writedata                       => mm_interconnect_0_flash_flash_erase_control_writedata,                   --                                                    .writedata
			Flash_flash_erase_control_byteenable                      => mm_interconnect_0_flash_flash_erase_control_byteenable,                  --                                                    .byteenable
			Flash_flash_erase_control_waitrequest                     => mm_interconnect_0_flash_flash_erase_control_waitrequest,                 --                                                    .waitrequest
			Flash_flash_erase_control_chipselect                      => mm_interconnect_0_flash_flash_erase_control_chipselect,                  --                                                    .chipselect
			Green_LEDs_avalon_parallel_port_slave_address             => mm_interconnect_0_green_leds_avalon_parallel_port_slave_address,         --               Green_LEDs_avalon_parallel_port_slave.address
			Green_LEDs_avalon_parallel_port_slave_write               => mm_interconnect_0_green_leds_avalon_parallel_port_slave_write,           --                                                    .write
			Green_LEDs_avalon_parallel_port_slave_read                => mm_interconnect_0_green_leds_avalon_parallel_port_slave_read,            --                                                    .read
			Green_LEDs_avalon_parallel_port_slave_readdata            => mm_interconnect_0_green_leds_avalon_parallel_port_slave_readdata,        --                                                    .readdata
			Green_LEDs_avalon_parallel_port_slave_writedata           => mm_interconnect_0_green_leds_avalon_parallel_port_slave_writedata,       --                                                    .writedata
			Green_LEDs_avalon_parallel_port_slave_byteenable          => mm_interconnect_0_green_leds_avalon_parallel_port_slave_byteenable,      --                                                    .byteenable
			Green_LEDs_avalon_parallel_port_slave_chipselect          => mm_interconnect_0_green_leds_avalon_parallel_port_slave_chipselect,      --                                                    .chipselect
			Interval_Timer_s1_address                                 => mm_interconnect_0_interval_timer_s1_address,                             --                                   Interval_Timer_s1.address
			Interval_Timer_s1_write                                   => mm_interconnect_0_interval_timer_s1_write,                               --                                                    .write
			Interval_Timer_s1_readdata                                => mm_interconnect_0_interval_timer_s1_readdata,                            --                                                    .readdata
			Interval_Timer_s1_writedata                               => mm_interconnect_0_interval_timer_s1_writedata,                           --                                                    .writedata
			Interval_Timer_s1_chipselect                              => mm_interconnect_0_interval_timer_s1_chipselect,                          --                                                    .chipselect
			JTAG_UART_avalon_jtag_slave_address                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,                   --                         JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write                         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                     --                                                    .write
			JTAG_UART_avalon_jtag_slave_read                          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                      --                                                    .read
			JTAG_UART_avalon_jtag_slave_readdata                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,                  --                                                    .readdata
			JTAG_UART_avalon_jtag_slave_writedata                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,                 --                                                    .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,               --                                                    .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,                --                                                    .chipselect
			JTAG_UART_2nd_Core_avalon_jtag_slave_address              => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address,          --                JTAG_UART_2nd_Core_avalon_jtag_slave.address
			JTAG_UART_2nd_Core_avalon_jtag_slave_write                => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write,            --                                                    .write
			JTAG_UART_2nd_Core_avalon_jtag_slave_read                 => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read,             --                                                    .read
			JTAG_UART_2nd_Core_avalon_jtag_slave_readdata             => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata,         --                                                    .readdata
			JTAG_UART_2nd_Core_avalon_jtag_slave_writedata            => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata,        --                                                    .writedata
			JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest          => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest,      --                                                    .waitrequest
			JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect           => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect,       --                                                    .chipselect
			Processor1_debug_mem_slave_address                        => mm_interconnect_0_processor1_debug_mem_slave_address,                    --                          Processor1_debug_mem_slave.address
			Processor1_debug_mem_slave_write                          => mm_interconnect_0_processor1_debug_mem_slave_write,                      --                                                    .write
			Processor1_debug_mem_slave_read                           => mm_interconnect_0_processor1_debug_mem_slave_read,                       --                                                    .read
			Processor1_debug_mem_slave_readdata                       => mm_interconnect_0_processor1_debug_mem_slave_readdata,                   --                                                    .readdata
			Processor1_debug_mem_slave_writedata                      => mm_interconnect_0_processor1_debug_mem_slave_writedata,                  --                                                    .writedata
			Processor1_debug_mem_slave_byteenable                     => mm_interconnect_0_processor1_debug_mem_slave_byteenable,                 --                                                    .byteenable
			Processor1_debug_mem_slave_waitrequest                    => mm_interconnect_0_processor1_debug_mem_slave_waitrequest,                --                                                    .waitrequest
			Processor1_debug_mem_slave_debugaccess                    => mm_interconnect_0_processor1_debug_mem_slave_debugaccess,                --                                                    .debugaccess
			Processor2_debug_mem_slave_address                        => mm_interconnect_0_processor2_debug_mem_slave_address,                    --                          Processor2_debug_mem_slave.address
			Processor2_debug_mem_slave_write                          => mm_interconnect_0_processor2_debug_mem_slave_write,                      --                                                    .write
			Processor2_debug_mem_slave_read                           => mm_interconnect_0_processor2_debug_mem_slave_read,                       --                                                    .read
			Processor2_debug_mem_slave_readdata                       => mm_interconnect_0_processor2_debug_mem_slave_readdata,                   --                                                    .readdata
			Processor2_debug_mem_slave_writedata                      => mm_interconnect_0_processor2_debug_mem_slave_writedata,                  --                                                    .writedata
			Processor2_debug_mem_slave_byteenable                     => mm_interconnect_0_processor2_debug_mem_slave_byteenable,                 --                                                    .byteenable
			Processor2_debug_mem_slave_waitrequest                    => mm_interconnect_0_processor2_debug_mem_slave_waitrequest,                --                                                    .waitrequest
			Processor2_debug_mem_slave_debugaccess                    => mm_interconnect_0_processor2_debug_mem_slave_debugaccess,                --                                                    .debugaccess
			Pushbuttons_avalon_parallel_port_slave_address            => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address,        --              Pushbuttons_avalon_parallel_port_slave.address
			Pushbuttons_avalon_parallel_port_slave_write              => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write,          --                                                    .write
			Pushbuttons_avalon_parallel_port_slave_read               => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read,           --                                                    .read
			Pushbuttons_avalon_parallel_port_slave_readdata           => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata,       --                                                    .readdata
			Pushbuttons_avalon_parallel_port_slave_writedata          => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata,      --                                                    .writedata
			Pushbuttons_avalon_parallel_port_slave_byteenable         => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable,     --                                                    .byteenable
			Pushbuttons_avalon_parallel_port_slave_chipselect         => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect,     --                                                    .chipselect
			Red_LEDs_avalon_parallel_port_slave_address               => mm_interconnect_0_red_leds_avalon_parallel_port_slave_address,           --                 Red_LEDs_avalon_parallel_port_slave.address
			Red_LEDs_avalon_parallel_port_slave_write                 => mm_interconnect_0_red_leds_avalon_parallel_port_slave_write,             --                                                    .write
			Red_LEDs_avalon_parallel_port_slave_read                  => mm_interconnect_0_red_leds_avalon_parallel_port_slave_read,              --                                                    .read
			Red_LEDs_avalon_parallel_port_slave_readdata              => mm_interconnect_0_red_leds_avalon_parallel_port_slave_readdata,          --                                                    .readdata
			Red_LEDs_avalon_parallel_port_slave_writedata             => mm_interconnect_0_red_leds_avalon_parallel_port_slave_writedata,         --                                                    .writedata
			Red_LEDs_avalon_parallel_port_slave_byteenable            => mm_interconnect_0_red_leds_avalon_parallel_port_slave_byteenable,        --                                                    .byteenable
			Red_LEDs_avalon_parallel_port_slave_chipselect            => mm_interconnect_0_red_leds_avalon_parallel_port_slave_chipselect,        --                                                    .chipselect
			SDRAM_s1_address                                          => mm_interconnect_0_sdram_s1_address,                                      --                                            SDRAM_s1.address
			SDRAM_s1_write                                            => mm_interconnect_0_sdram_s1_write,                                        --                                                    .write
			SDRAM_s1_read                                             => mm_interconnect_0_sdram_s1_read,                                         --                                                    .read
			SDRAM_s1_readdata                                         => mm_interconnect_0_sdram_s1_readdata,                                     --                                                    .readdata
			SDRAM_s1_writedata                                        => mm_interconnect_0_sdram_s1_writedata,                                    --                                                    .writedata
			SDRAM_s1_byteenable                                       => mm_interconnect_0_sdram_s1_byteenable,                                   --                                                    .byteenable
			SDRAM_s1_readdatavalid                                    => mm_interconnect_0_sdram_s1_readdatavalid,                                --                                                    .readdatavalid
			SDRAM_s1_waitrequest                                      => mm_interconnect_0_sdram_s1_waitrequest,                                  --                                                    .waitrequest
			SDRAM_s1_chipselect                                       => mm_interconnect_0_sdram_s1_chipselect,                                   --                                                    .chipselect
			Serial_Port_avalon_rs232_slave_address                    => mm_interconnect_0_serial_port_avalon_rs232_slave_address,                --                      Serial_Port_avalon_rs232_slave.address
			Serial_Port_avalon_rs232_slave_write                      => mm_interconnect_0_serial_port_avalon_rs232_slave_write,                  --                                                    .write
			Serial_Port_avalon_rs232_slave_read                       => mm_interconnect_0_serial_port_avalon_rs232_slave_read,                   --                                                    .read
			Serial_Port_avalon_rs232_slave_readdata                   => mm_interconnect_0_serial_port_avalon_rs232_slave_readdata,               --                                                    .readdata
			Serial_Port_avalon_rs232_slave_writedata                  => mm_interconnect_0_serial_port_avalon_rs232_slave_writedata,              --                                                    .writedata
			Serial_Port_avalon_rs232_slave_byteenable                 => mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable,             --                                                    .byteenable
			Serial_Port_avalon_rs232_slave_chipselect                 => mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect,             --                                                    .chipselect
			Slider_Switches_avalon_parallel_port_slave_address        => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_address,    --          Slider_Switches_avalon_parallel_port_slave.address
			Slider_Switches_avalon_parallel_port_slave_write          => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_write,      --                                                    .write
			Slider_Switches_avalon_parallel_port_slave_read           => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_read,       --                                                    .read
			Slider_Switches_avalon_parallel_port_slave_readdata       => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_readdata,   --                                                    .readdata
			Slider_Switches_avalon_parallel_port_slave_writedata      => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_writedata,  --                                                    .writedata
			Slider_Switches_avalon_parallel_port_slave_byteenable     => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_byteenable, --                                                    .byteenable
			Slider_Switches_avalon_parallel_port_slave_chipselect     => mm_interconnect_0_slider_switches_avalon_parallel_port_slave_chipselect, --                                                    .chipselect
			SRAM_avalon_sram_slave_address                            => mm_interconnect_0_sram_avalon_sram_slave_address,                        --                              SRAM_avalon_sram_slave.address
			SRAM_avalon_sram_slave_write                              => mm_interconnect_0_sram_avalon_sram_slave_write,                          --                                                    .write
			SRAM_avalon_sram_slave_read                               => mm_interconnect_0_sram_avalon_sram_slave_read,                           --                                                    .read
			SRAM_avalon_sram_slave_readdata                           => mm_interconnect_0_sram_avalon_sram_slave_readdata,                       --                                                    .readdata
			SRAM_avalon_sram_slave_writedata                          => mm_interconnect_0_sram_avalon_sram_slave_writedata,                      --                                                    .writedata
			SRAM_avalon_sram_slave_byteenable                         => mm_interconnect_0_sram_avalon_sram_slave_byteenable,                     --                                                    .byteenable
			SRAM_avalon_sram_slave_readdatavalid                      => mm_interconnect_0_sram_avalon_sram_slave_readdatavalid,                  --                                                    .readdatavalid
			SysID_control_slave_address                               => mm_interconnect_0_sysid_control_slave_address,                           --                                 SysID_control_slave.address
			SysID_control_slave_readdata                              => mm_interconnect_0_sysid_control_slave_readdata                           --                                                    .readdata
		);

	irq_mapper : component nios_system_irq_mapper
		port map (
			clk           => system_pll_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			sender_irq    => processor1_irq_irq                  --    sender.irq
		);

	irq_mapper_001 : component nios_system_irq_mapper
		port map (
			clk           => system_pll_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_001_receiver5_irq,       -- receiver5.irq
			sender_irq    => processor2_irq_irq                  --    sender.irq
		);

	rst_controller : component nios_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => system_pll_reset_source_reset,  -- reset_in0.reset
			clk            => system_pll_sys_clk_clk,         --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component nios_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => processor1_debug_reset_request_reset,   -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,          -- reset_in1.reset
			clk            => system_pll_sys_clk_clk,                 --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component nios_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => processor2_debug_reset_request_reset,   -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,          -- reset_in1.reset
			clk            => system_pll_sys_clk_clk,                 --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	system_pll_reset_source_reset_ports_inv <= not system_pll_reset_source_reset;

	mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write;

	mm_interconnect_0_interval_timer_s1_write_ports_inv <= not mm_interconnect_0_interval_timer_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of nios_system
