-- nios_system_Video_In_Subsystem_Edge_Detection_Subsystem.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_system_Video_In_Subsystem_Edge_Detection_Subsystem is
	port (
		edge_detection_control_slave_address    : in  std_logic_vector(1 downto 0)  := (others => '0'); -- edge_detection_control_slave.address
		edge_detection_control_slave_write_n    : in  std_logic                     := '0';             --                             .write_n
		edge_detection_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                             .writedata
		edge_detection_control_slave_chipselect : in  std_logic                     := '0';             --                             .chipselect
		edge_detection_control_slave_readdata   : out std_logic_vector(31 downto 0);                    --                             .readdata
		sys_clk_clk                             : in  std_logic                     := '0';             --                      sys_clk.clk
		sys_reset_reset_n                       : in  std_logic                     := '0';             --                    sys_reset.reset_n
		video_stream_sink_data                  : in  std_logic_vector(23 downto 0) := (others => '0'); --            video_stream_sink.data
		video_stream_sink_startofpacket         : in  std_logic                     := '0';             --                             .startofpacket
		video_stream_sink_endofpacket           : in  std_logic                     := '0';             --                             .endofpacket
		video_stream_sink_valid                 : in  std_logic                     := '0';             --                             .valid
		video_stream_sink_ready                 : out std_logic;                                        --                             .ready
		video_stream_source_ready               : in  std_logic                     := '0';             --          video_stream_source.ready
		video_stream_source_data                : out std_logic_vector(23 downto 0);                    --                             .data
		video_stream_source_startofpacket       : out std_logic;                                        --                             .startofpacket
		video_stream_source_endofpacket         : out std_logic;                                        --                             .endofpacket
		video_stream_source_valid               : out std_logic                                         --                             .valid
	);
end entity nios_system_Video_In_Subsystem_Edge_Detection_Subsystem;

architecture rtl of nios_system_Video_In_Subsystem_Edge_Detection_Subsystem is
	component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Chroma_Filter is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(7 downto 0)                      -- data
		);
	end component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Chroma_Filter;

	component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Chroma_Upsampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(23 downto 0)                     -- data
		);
	end component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Chroma_Upsampler;

	component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Edge_Detection is
		port (
			clk               : in  std_logic                    := 'X';             -- clk
			reset             : in  std_logic                    := 'X';             -- reset
			in_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			in_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			in_valid          : in  std_logic                    := 'X';             -- valid
			in_ready          : out std_logic;                                       -- ready
			out_ready         : in  std_logic                    := 'X';             -- ready
			out_data          : out std_logic_vector(7 downto 0);                    -- data
			out_startofpacket : out std_logic;                                       -- startofpacket
			out_endofpacket   : out std_logic;                                       -- endofpacket
			out_valid         : out std_logic                                        -- valid
		);
	end component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Edge_Detection;

	component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Edge_Detection_Router_Controller is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Edge_Detection_Router_Controller;

	component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Video_Stream_Merger is
		port (
			clk                       : in  std_logic                     := 'X';             -- clk
			reset                     : in  std_logic                     := 'X';             -- reset
			stream_in_data_0          : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket_0 : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket_0   : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid_0         : in  std_logic                     := 'X';             -- valid
			stream_in_ready_0         : out std_logic;                                        -- ready
			stream_in_data_1          : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket_1 : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket_1   : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid_1         : in  std_logic                     := 'X';             -- valid
			stream_in_ready_1         : out std_logic;                                        -- ready
			sync_data                 : in  std_logic                     := 'X';             -- data
			sync_valid                : in  std_logic                     := 'X';             -- valid
			sync_ready                : out std_logic;                                        -- ready
			stream_out_ready          : in  std_logic                     := 'X';             -- ready
			stream_out_data           : out std_logic_vector(23 downto 0);                    -- data
			stream_out_startofpacket  : out std_logic;                                        -- startofpacket
			stream_out_endofpacket    : out std_logic;                                        -- endofpacket
			stream_out_valid          : out std_logic                                         -- valid
		);
	end component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Video_Stream_Merger;

	component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Video_Stream_Splitter is
		port (
			clk                        : in  std_logic                     := 'X';             -- clk
			reset                      : in  std_logic                     := 'X';             -- reset
			stream_in_data             : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket    : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket      : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid            : in  std_logic                     := 'X';             -- valid
			stream_in_ready            : out std_logic;                                        -- ready
			sync_ready                 : in  std_logic                     := 'X';             -- ready
			sync_data                  : out std_logic;                                        -- data
			sync_valid                 : out std_logic;                                        -- valid
			stream_out_ready_0         : in  std_logic                     := 'X';             -- ready
			stream_out_data_0          : out std_logic_vector(23 downto 0);                    -- data
			stream_out_startofpacket_0 : out std_logic;                                        -- startofpacket
			stream_out_endofpacket_0   : out std_logic;                                        -- endofpacket
			stream_out_valid_0         : out std_logic;                                        -- valid
			stream_out_ready_1         : in  std_logic                     := 'X';             -- ready
			stream_out_data_1          : out std_logic_vector(23 downto 0);                    -- data
			stream_out_startofpacket_1 : out std_logic;                                        -- startofpacket
			stream_out_endofpacket_1   : out std_logic;                                        -- endofpacket
			stream_out_valid_1         : out std_logic;                                        -- valid
			stream_select              : in  std_logic                     := 'X'              -- export
		);
	end component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Video_Stream_Splitter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal chroma_filter_avalon_chroma_source_valid                          : std_logic;                     -- Chroma_Filter:stream_out_valid -> Edge_Detection:in_valid
	signal chroma_filter_avalon_chroma_source_data                           : std_logic_vector(7 downto 0);  -- Chroma_Filter:stream_out_data -> Edge_Detection:in_data
	signal chroma_filter_avalon_chroma_source_ready                          : std_logic;                     -- Edge_Detection:in_ready -> Chroma_Filter:stream_out_ready
	signal chroma_filter_avalon_chroma_source_startofpacket                  : std_logic;                     -- Chroma_Filter:stream_out_startofpacket -> Edge_Detection:in_startofpacket
	signal chroma_filter_avalon_chroma_source_endofpacket                    : std_logic;                     -- Chroma_Filter:stream_out_endofpacket -> Edge_Detection:in_endofpacket
	signal chroma_upsampler_avalon_chroma_source_valid                       : std_logic;                     -- Chroma_Upsampler:stream_out_valid -> Video_Stream_Merger:stream_in_valid_1
	signal chroma_upsampler_avalon_chroma_source_data                        : std_logic_vector(23 downto 0); -- Chroma_Upsampler:stream_out_data -> Video_Stream_Merger:stream_in_data_1
	signal chroma_upsampler_avalon_chroma_source_ready                       : std_logic;                     -- Video_Stream_Merger:stream_in_ready_1 -> Chroma_Upsampler:stream_out_ready
	signal chroma_upsampler_avalon_chroma_source_startofpacket               : std_logic;                     -- Chroma_Upsampler:stream_out_startofpacket -> Video_Stream_Merger:stream_in_startofpacket_1
	signal chroma_upsampler_avalon_chroma_source_endofpacket                 : std_logic;                     -- Chroma_Upsampler:stream_out_endofpacket -> Video_Stream_Merger:stream_in_endofpacket_1
	signal edge_detection_avalon_edge_detection_source_valid                 : std_logic;                     -- Edge_Detection:out_valid -> Chroma_Upsampler:stream_in_valid
	signal edge_detection_avalon_edge_detection_source_data                  : std_logic_vector(7 downto 0);  -- Edge_Detection:out_data -> Chroma_Upsampler:stream_in_data
	signal edge_detection_avalon_edge_detection_source_ready                 : std_logic;                     -- Chroma_Upsampler:stream_in_ready -> Edge_Detection:out_ready
	signal edge_detection_avalon_edge_detection_source_startofpacket         : std_logic;                     -- Edge_Detection:out_startofpacket -> Chroma_Upsampler:stream_in_startofpacket
	signal edge_detection_avalon_edge_detection_source_endofpacket           : std_logic;                     -- Edge_Detection:out_endofpacket -> Chroma_Upsampler:stream_in_endofpacket
	signal video_stream_splitter_avalon_stream_router_source_0_valid         : std_logic;                     -- Video_Stream_Splitter:stream_out_valid_0 -> Video_Stream_Merger:stream_in_valid_0
	signal video_stream_splitter_avalon_stream_router_source_0_data          : std_logic_vector(23 downto 0); -- Video_Stream_Splitter:stream_out_data_0 -> Video_Stream_Merger:stream_in_data_0
	signal video_stream_splitter_avalon_stream_router_source_0_ready         : std_logic;                     -- Video_Stream_Merger:stream_in_ready_0 -> Video_Stream_Splitter:stream_out_ready_0
	signal video_stream_splitter_avalon_stream_router_source_0_startofpacket : std_logic;                     -- Video_Stream_Splitter:stream_out_startofpacket_0 -> Video_Stream_Merger:stream_in_startofpacket_0
	signal video_stream_splitter_avalon_stream_router_source_0_endofpacket   : std_logic;                     -- Video_Stream_Splitter:stream_out_endofpacket_0 -> Video_Stream_Merger:stream_in_endofpacket_0
	signal video_stream_splitter_avalon_stream_router_source_1_valid         : std_logic;                     -- Video_Stream_Splitter:stream_out_valid_1 -> Chroma_Filter:stream_in_valid
	signal video_stream_splitter_avalon_stream_router_source_1_data          : std_logic_vector(23 downto 0); -- Video_Stream_Splitter:stream_out_data_1 -> Chroma_Filter:stream_in_data
	signal video_stream_splitter_avalon_stream_router_source_1_ready         : std_logic;                     -- Chroma_Filter:stream_in_ready -> Video_Stream_Splitter:stream_out_ready_1
	signal video_stream_splitter_avalon_stream_router_source_1_startofpacket : std_logic;                     -- Video_Stream_Splitter:stream_out_startofpacket_1 -> Chroma_Filter:stream_in_startofpacket
	signal video_stream_splitter_avalon_stream_router_source_1_endofpacket   : std_logic;                     -- Video_Stream_Splitter:stream_out_endofpacket_1 -> Chroma_Filter:stream_in_endofpacket
	signal video_stream_splitter_avalon_sync_source_valid                    : std_logic;                     -- Video_Stream_Splitter:sync_valid -> Video_Stream_Merger:sync_valid
	signal video_stream_splitter_avalon_sync_source_data                     : std_logic;                     -- Video_Stream_Splitter:sync_data -> Video_Stream_Merger:sync_data
	signal video_stream_splitter_avalon_sync_source_ready                    : std_logic;                     -- Video_Stream_Merger:sync_ready -> Video_Stream_Splitter:sync_ready
	signal edge_detection_router_controller_external_connection_export       : std_logic;                     -- Edge_Detection_Router_Controller:out_port -> Video_Stream_Splitter:stream_select
	signal rst_controller_reset_out_reset                                    : std_logic;                     -- rst_controller:reset_out -> [Chroma_Filter:reset, Chroma_Upsampler:reset, Edge_Detection:reset, Video_Stream_Merger:reset, Video_Stream_Splitter:reset, rst_controller_reset_out_reset:in]
	signal sys_reset_reset_n_ports_inv                                       : std_logic;                     -- sys_reset_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv                          : std_logic;                     -- rst_controller_reset_out_reset:inv -> Edge_Detection_Router_Controller:reset_n

begin

	chroma_filter : component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Chroma_Filter
		port map (
			clk                      => sys_clk_clk,                                                       --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                                    --                reset.reset
			stream_in_startofpacket  => video_stream_splitter_avalon_stream_router_source_1_startofpacket, --   avalon_chroma_sink.startofpacket
			stream_in_endofpacket    => video_stream_splitter_avalon_stream_router_source_1_endofpacket,   --                     .endofpacket
			stream_in_valid          => video_stream_splitter_avalon_stream_router_source_1_valid,         --                     .valid
			stream_in_ready          => video_stream_splitter_avalon_stream_router_source_1_ready,         --                     .ready
			stream_in_data           => video_stream_splitter_avalon_stream_router_source_1_data,          --                     .data
			stream_out_ready         => chroma_filter_avalon_chroma_source_ready,                          -- avalon_chroma_source.ready
			stream_out_startofpacket => chroma_filter_avalon_chroma_source_startofpacket,                  --                     .startofpacket
			stream_out_endofpacket   => chroma_filter_avalon_chroma_source_endofpacket,                    --                     .endofpacket
			stream_out_valid         => chroma_filter_avalon_chroma_source_valid,                          --                     .valid
			stream_out_data          => chroma_filter_avalon_chroma_source_data                            --                     .data
		);

	chroma_upsampler : component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Chroma_Upsampler
		port map (
			clk                      => sys_clk_clk,                                               --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                            --                reset.reset
			stream_in_startofpacket  => edge_detection_avalon_edge_detection_source_startofpacket, --   avalon_chroma_sink.startofpacket
			stream_in_endofpacket    => edge_detection_avalon_edge_detection_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => edge_detection_avalon_edge_detection_source_valid,         --                     .valid
			stream_in_ready          => edge_detection_avalon_edge_detection_source_ready,         --                     .ready
			stream_in_data           => edge_detection_avalon_edge_detection_source_data,          --                     .data
			stream_out_ready         => chroma_upsampler_avalon_chroma_source_ready,               -- avalon_chroma_source.ready
			stream_out_startofpacket => chroma_upsampler_avalon_chroma_source_startofpacket,       --                     .startofpacket
			stream_out_endofpacket   => chroma_upsampler_avalon_chroma_source_endofpacket,         --                     .endofpacket
			stream_out_valid         => chroma_upsampler_avalon_chroma_source_valid,               --                     .valid
			stream_out_data          => chroma_upsampler_avalon_chroma_source_data                 --                     .data
		);

	edge_detection : component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Edge_Detection
		port map (
			clk               => sys_clk_clk,                                               --                          clk.clk
			reset             => rst_controller_reset_out_reset,                            --                        reset.reset
			in_data           => chroma_filter_avalon_chroma_source_data,                   --   avalon_edge_detection_sink.data
			in_startofpacket  => chroma_filter_avalon_chroma_source_startofpacket,          --                             .startofpacket
			in_endofpacket    => chroma_filter_avalon_chroma_source_endofpacket,            --                             .endofpacket
			in_valid          => chroma_filter_avalon_chroma_source_valid,                  --                             .valid
			in_ready          => chroma_filter_avalon_chroma_source_ready,                  --                             .ready
			out_ready         => edge_detection_avalon_edge_detection_source_ready,         -- avalon_edge_detection_source.ready
			out_data          => edge_detection_avalon_edge_detection_source_data,          --                             .data
			out_startofpacket => edge_detection_avalon_edge_detection_source_startofpacket, --                             .startofpacket
			out_endofpacket   => edge_detection_avalon_edge_detection_source_endofpacket,   --                             .endofpacket
			out_valid         => edge_detection_avalon_edge_detection_source_valid          --                             .valid
		);

	edge_detection_router_controller : component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Edge_Detection_Router_Controller
		port map (
			clk        => sys_clk_clk,                                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                    --               reset.reset_n
			address    => edge_detection_control_slave_address,                        --                  s1.address
			write_n    => edge_detection_control_slave_write_n,                        --                    .write_n
			writedata  => edge_detection_control_slave_writedata,                      --                    .writedata
			chipselect => edge_detection_control_slave_chipselect,                     --                    .chipselect
			readdata   => edge_detection_control_slave_readdata,                       --                    .readdata
			out_port   => edge_detection_router_controller_external_connection_export  -- external_connection.export
		);

	video_stream_merger : component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Video_Stream_Merger
		port map (
			clk                       => sys_clk_clk,                                                       --                         clk.clk
			reset                     => rst_controller_reset_out_reset,                                    --                       reset.reset
			stream_in_data_0          => video_stream_splitter_avalon_stream_router_source_0_data,          -- avalon_stream_router_sink_0.data
			stream_in_startofpacket_0 => video_stream_splitter_avalon_stream_router_source_0_startofpacket, --                            .startofpacket
			stream_in_endofpacket_0   => video_stream_splitter_avalon_stream_router_source_0_endofpacket,   --                            .endofpacket
			stream_in_valid_0         => video_stream_splitter_avalon_stream_router_source_0_valid,         --                            .valid
			stream_in_ready_0         => video_stream_splitter_avalon_stream_router_source_0_ready,         --                            .ready
			stream_in_data_1          => chroma_upsampler_avalon_chroma_source_data,                        -- avalon_stream_router_sink_1.data
			stream_in_startofpacket_1 => chroma_upsampler_avalon_chroma_source_startofpacket,               --                            .startofpacket
			stream_in_endofpacket_1   => chroma_upsampler_avalon_chroma_source_endofpacket,                 --                            .endofpacket
			stream_in_valid_1         => chroma_upsampler_avalon_chroma_source_valid,                       --                            .valid
			stream_in_ready_1         => chroma_upsampler_avalon_chroma_source_ready,                       --                            .ready
			sync_data                 => video_stream_splitter_avalon_sync_source_data,                     --            avalon_sync_sink.data
			sync_valid                => video_stream_splitter_avalon_sync_source_valid,                    --                            .valid
			sync_ready                => video_stream_splitter_avalon_sync_source_ready,                    --                            .ready
			stream_out_ready          => video_stream_source_ready,                                         -- avalon_stream_router_source.ready
			stream_out_data           => video_stream_source_data,                                          --                            .data
			stream_out_startofpacket  => video_stream_source_startofpacket,                                 --                            .startofpacket
			stream_out_endofpacket    => video_stream_source_endofpacket,                                   --                            .endofpacket
			stream_out_valid          => video_stream_source_valid                                          --                            .valid
		);

	video_stream_splitter : component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem_Video_Stream_Splitter
		port map (
			clk                        => sys_clk_clk,                                                       --                           clk.clk
			reset                      => rst_controller_reset_out_reset,                                    --                         reset.reset
			stream_in_data             => video_stream_sink_data,                                            --     avalon_stream_router_sink.data
			stream_in_startofpacket    => video_stream_sink_startofpacket,                                   --                              .startofpacket
			stream_in_endofpacket      => video_stream_sink_endofpacket,                                     --                              .endofpacket
			stream_in_valid            => video_stream_sink_valid,                                           --                              .valid
			stream_in_ready            => video_stream_sink_ready,                                           --                              .ready
			sync_ready                 => video_stream_splitter_avalon_sync_source_ready,                    --            avalon_sync_source.ready
			sync_data                  => video_stream_splitter_avalon_sync_source_data,                     --                              .data
			sync_valid                 => video_stream_splitter_avalon_sync_source_valid,                    --                              .valid
			stream_out_ready_0         => video_stream_splitter_avalon_stream_router_source_0_ready,         -- avalon_stream_router_source_0.ready
			stream_out_data_0          => video_stream_splitter_avalon_stream_router_source_0_data,          --                              .data
			stream_out_startofpacket_0 => video_stream_splitter_avalon_stream_router_source_0_startofpacket, --                              .startofpacket
			stream_out_endofpacket_0   => video_stream_splitter_avalon_stream_router_source_0_endofpacket,   --                              .endofpacket
			stream_out_valid_0         => video_stream_splitter_avalon_stream_router_source_0_valid,         --                              .valid
			stream_out_ready_1         => video_stream_splitter_avalon_stream_router_source_1_ready,         -- avalon_stream_router_source_1.ready
			stream_out_data_1          => video_stream_splitter_avalon_stream_router_source_1_data,          --                              .data
			stream_out_startofpacket_1 => video_stream_splitter_avalon_stream_router_source_1_startofpacket, --                              .startofpacket
			stream_out_endofpacket_1   => video_stream_splitter_avalon_stream_router_source_1_endofpacket,   --                              .endofpacket
			stream_out_valid_1         => video_stream_splitter_avalon_stream_router_source_1_valid,         --                              .valid
			stream_select              => edge_detection_router_controller_external_connection_export        --            external_interface.export
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_reset_reset_n_ports_inv,    -- reset_in0.reset
			clk            => sys_clk_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	sys_reset_reset_n_ports_inv <= not sys_reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_system_Video_In_Subsystem_Edge_Detection_Subsystem
