-- nios_system_Video_In_Subsystem.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_system_Video_In_Subsystem is
	port (
		edge_detection_control_slave_address    : in  std_logic_vector(1 downto 0)  := (others => '0'); -- edge_detection_control_slave.address
		edge_detection_control_slave_write_n    : in  std_logic                     := '0';             --                             .write_n
		edge_detection_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                             .writedata
		edge_detection_control_slave_chipselect : in  std_logic                     := '0';             --                             .chipselect
		edge_detection_control_slave_readdata   : out std_logic_vector(31 downto 0);                    --                             .readdata
		sys_clk_clk                             : in  std_logic                     := '0';             --                      sys_clk.clk
		sys_reset_reset_n                       : in  std_logic                     := '0';             --                    sys_reset.reset_n
		video_in_TD_CLK27                       : in  std_logic                     := '0';             --                     video_in.TD_CLK27
		video_in_TD_DATA                        : in  std_logic_vector(7 downto 0)  := (others => '0'); --                             .TD_DATA
		video_in_TD_HS                          : in  std_logic                     := '0';             --                             .TD_HS
		video_in_TD_VS                          : in  std_logic                     := '0';             --                             .TD_VS
		video_in_clk27_reset                    : in  std_logic                     := '0';             --                             .clk27_reset
		video_in_TD_RESET                       : out std_logic;                                        --                             .TD_RESET
		video_in_overflow_flag                  : out std_logic;                                        --                             .overflow_flag
		video_in_dma_control_slave_address      : in  std_logic_vector(1 downto 0)  := (others => '0'); --   video_in_dma_control_slave.address
		video_in_dma_control_slave_byteenable   : in  std_logic_vector(3 downto 0)  := (others => '0'); --                             .byteenable
		video_in_dma_control_slave_read         : in  std_logic                     := '0';             --                             .read
		video_in_dma_control_slave_write        : in  std_logic                     := '0';             --                             .write
		video_in_dma_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => '0'); --                             .writedata
		video_in_dma_control_slave_readdata     : out std_logic_vector(31 downto 0);                    --                             .readdata
		video_in_dma_master_address             : out std_logic_vector(31 downto 0);                    --          video_in_dma_master.address
		video_in_dma_master_waitrequest         : in  std_logic                     := '0';             --                             .waitrequest
		video_in_dma_master_write               : out std_logic;                                        --                             .write
		video_in_dma_master_writedata           : out std_logic_vector(15 downto 0)                     --                             .writedata
	);
end entity nios_system_Video_In_Subsystem;

architecture rtl of nios_system_Video_In_Subsystem is
	component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem is
		port (
			edge_detection_control_slave_address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			edge_detection_control_slave_write_n    : in  std_logic                     := 'X';             -- write_n
			edge_detection_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			edge_detection_control_slave_chipselect : in  std_logic                     := 'X';             -- chipselect
			edge_detection_control_slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			sys_clk_clk                             : in  std_logic                     := 'X';             -- clk
			sys_reset_reset_n                       : in  std_logic                     := 'X';             -- reset_n
			video_stream_sink_data                  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			video_stream_sink_startofpacket         : in  std_logic                     := 'X';             -- startofpacket
			video_stream_sink_endofpacket           : in  std_logic                     := 'X';             -- endofpacket
			video_stream_sink_valid                 : in  std_logic                     := 'X';             -- valid
			video_stream_sink_ready                 : out std_logic;                                        -- ready
			video_stream_source_ready               : in  std_logic                     := 'X';             -- ready
			video_stream_source_data                : out std_logic_vector(23 downto 0);                    -- data
			video_stream_source_startofpacket       : out std_logic;                                        -- startofpacket
			video_stream_source_endofpacket         : out std_logic;                                        -- endofpacket
			video_stream_source_valid               : out std_logic                                         -- valid
		);
	end component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem;

	component nios_system_Video_In_Subsystem_Video_In is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(15 downto 0);                    -- data
			TD_CLK27                 : in  std_logic                     := 'X';             -- export
			TD_DATA                  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			TD_HS                    : in  std_logic                     := 'X';             -- export
			TD_VS                    : in  std_logic                     := 'X';             -- export
			clk27_reset              : in  std_logic                     := 'X';             -- export
			TD_RESET                 : out std_logic;                                        -- export
			overflow_flag            : out std_logic                                         -- export
		);
	end component nios_system_Video_In_Subsystem_Video_In;

	component nios_system_Video_In_Subsystem_Video_In_CSC is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(23 downto 0)                     -- data
		);
	end component nios_system_Video_In_Subsystem_Video_In_CSC;

	component nios_system_Video_In_Subsystem_Video_In_Chroma_Resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(23 downto 0)                     -- data
		);
	end component nios_system_Video_In_Subsystem_Video_In_Chroma_Resampler;

	component nios_system_Video_In_Subsystem_Video_In_Clipper is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_data          : out std_logic_vector(15 downto 0);                    -- data
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic                                         -- valid
		);
	end component nios_system_Video_In_Subsystem_Video_In_Clipper;

	component nios_system_Video_In_Subsystem_Video_In_DMA is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			stream_data          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			stream_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			stream_valid         : in  std_logic                     := 'X';             -- valid
			stream_ready         : out std_logic;                                        -- ready
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(15 downto 0)                     -- writedata
		);
	end component nios_system_Video_In_Subsystem_Video_In_DMA;

	component nios_system_Video_In_Subsystem_Video_In_RGB_Resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(15 downto 0)                     -- data
		);
	end component nios_system_Video_In_Subsystem_Video_In_RGB_Resampler;

	component nios_system_Video_In_Subsystem_Video_In_Scaler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(15 downto 0)                     -- data
		);
	end component nios_system_Video_In_Subsystem_Video_In_Scaler;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal video_in_chroma_resampler_avalon_chroma_source_valid         : std_logic;                     -- Video_In_Chroma_Resampler:stream_out_valid -> Edge_Detection_Subsystem:video_stream_sink_valid
	signal video_in_chroma_resampler_avalon_chroma_source_data          : std_logic_vector(23 downto 0); -- Video_In_Chroma_Resampler:stream_out_data -> Edge_Detection_Subsystem:video_stream_sink_data
	signal video_in_chroma_resampler_avalon_chroma_source_ready         : std_logic;                     -- Edge_Detection_Subsystem:video_stream_sink_ready -> Video_In_Chroma_Resampler:stream_out_ready
	signal video_in_chroma_resampler_avalon_chroma_source_startofpacket : std_logic;                     -- Video_In_Chroma_Resampler:stream_out_startofpacket -> Edge_Detection_Subsystem:video_stream_sink_startofpacket
	signal video_in_chroma_resampler_avalon_chroma_source_endofpacket   : std_logic;                     -- Video_In_Chroma_Resampler:stream_out_endofpacket -> Edge_Detection_Subsystem:video_stream_sink_endofpacket
	signal video_in_clipper_avalon_clipper_source_valid                 : std_logic;                     -- Video_In_Clipper:stream_out_valid -> Video_In_Scaler:stream_in_valid
	signal video_in_clipper_avalon_clipper_source_data                  : std_logic_vector(15 downto 0); -- Video_In_Clipper:stream_out_data -> Video_In_Scaler:stream_in_data
	signal video_in_clipper_avalon_clipper_source_ready                 : std_logic;                     -- Video_In_Scaler:stream_in_ready -> Video_In_Clipper:stream_out_ready
	signal video_in_clipper_avalon_clipper_source_startofpacket         : std_logic;                     -- Video_In_Clipper:stream_out_startofpacket -> Video_In_Scaler:stream_in_startofpacket
	signal video_in_clipper_avalon_clipper_source_endofpacket           : std_logic;                     -- Video_In_Clipper:stream_out_endofpacket -> Video_In_Scaler:stream_in_endofpacket
	signal video_in_csc_avalon_csc_source_valid                         : std_logic;                     -- Video_In_CSC:stream_out_valid -> Video_In_RGB_Resampler:stream_in_valid
	signal video_in_csc_avalon_csc_source_data                          : std_logic_vector(23 downto 0); -- Video_In_CSC:stream_out_data -> Video_In_RGB_Resampler:stream_in_data
	signal video_in_csc_avalon_csc_source_ready                         : std_logic;                     -- Video_In_RGB_Resampler:stream_in_ready -> Video_In_CSC:stream_out_ready
	signal video_in_csc_avalon_csc_source_startofpacket                 : std_logic;                     -- Video_In_CSC:stream_out_startofpacket -> Video_In_RGB_Resampler:stream_in_startofpacket
	signal video_in_csc_avalon_csc_source_endofpacket                   : std_logic;                     -- Video_In_CSC:stream_out_endofpacket -> Video_In_RGB_Resampler:stream_in_endofpacket
	signal video_in_avalon_decoder_source_valid                         : std_logic;                     -- Video_In:stream_out_valid -> Video_In_Chroma_Resampler:stream_in_valid
	signal video_in_avalon_decoder_source_data                          : std_logic_vector(15 downto 0); -- Video_In:stream_out_data -> Video_In_Chroma_Resampler:stream_in_data
	signal video_in_avalon_decoder_source_ready                         : std_logic;                     -- Video_In_Chroma_Resampler:stream_in_ready -> Video_In:stream_out_ready
	signal video_in_avalon_decoder_source_startofpacket                 : std_logic;                     -- Video_In:stream_out_startofpacket -> Video_In_Chroma_Resampler:stream_in_startofpacket
	signal video_in_avalon_decoder_source_endofpacket                   : std_logic;                     -- Video_In:stream_out_endofpacket -> Video_In_Chroma_Resampler:stream_in_endofpacket
	signal video_in_rgb_resampler_avalon_rgb_source_valid               : std_logic;                     -- Video_In_RGB_Resampler:stream_out_valid -> Video_In_Clipper:stream_in_valid
	signal video_in_rgb_resampler_avalon_rgb_source_data                : std_logic_vector(15 downto 0); -- Video_In_RGB_Resampler:stream_out_data -> Video_In_Clipper:stream_in_data
	signal video_in_rgb_resampler_avalon_rgb_source_ready               : std_logic;                     -- Video_In_Clipper:stream_in_ready -> Video_In_RGB_Resampler:stream_out_ready
	signal video_in_rgb_resampler_avalon_rgb_source_startofpacket       : std_logic;                     -- Video_In_RGB_Resampler:stream_out_startofpacket -> Video_In_Clipper:stream_in_startofpacket
	signal video_in_rgb_resampler_avalon_rgb_source_endofpacket         : std_logic;                     -- Video_In_RGB_Resampler:stream_out_endofpacket -> Video_In_Clipper:stream_in_endofpacket
	signal video_in_scaler_avalon_scaler_source_valid                   : std_logic;                     -- Video_In_Scaler:stream_out_valid -> Video_In_DMA:stream_valid
	signal video_in_scaler_avalon_scaler_source_data                    : std_logic_vector(15 downto 0); -- Video_In_Scaler:stream_out_data -> Video_In_DMA:stream_data
	signal video_in_scaler_avalon_scaler_source_ready                   : std_logic;                     -- Video_In_DMA:stream_ready -> Video_In_Scaler:stream_out_ready
	signal video_in_scaler_avalon_scaler_source_startofpacket           : std_logic;                     -- Video_In_Scaler:stream_out_startofpacket -> Video_In_DMA:stream_startofpacket
	signal video_in_scaler_avalon_scaler_source_endofpacket             : std_logic;                     -- Video_In_Scaler:stream_out_endofpacket -> Video_In_DMA:stream_endofpacket
	signal edge_detection_subsystem_video_stream_source_valid           : std_logic;                     -- Edge_Detection_Subsystem:video_stream_source_valid -> Video_In_CSC:stream_in_valid
	signal edge_detection_subsystem_video_stream_source_data            : std_logic_vector(23 downto 0); -- Edge_Detection_Subsystem:video_stream_source_data -> Video_In_CSC:stream_in_data
	signal edge_detection_subsystem_video_stream_source_ready           : std_logic;                     -- Video_In_CSC:stream_in_ready -> Edge_Detection_Subsystem:video_stream_source_ready
	signal edge_detection_subsystem_video_stream_source_startofpacket   : std_logic;                     -- Edge_Detection_Subsystem:video_stream_source_startofpacket -> Video_In_CSC:stream_in_startofpacket
	signal edge_detection_subsystem_video_stream_source_endofpacket     : std_logic;                     -- Edge_Detection_Subsystem:video_stream_source_endofpacket -> Video_In_CSC:stream_in_endofpacket
	signal rst_controller_reset_out_reset                               : std_logic;                     -- rst_controller:reset_out -> [Video_In:reset, Video_In_CSC:reset, Video_In_Chroma_Resampler:reset, Video_In_Clipper:reset, Video_In_DMA:reset, Video_In_RGB_Resampler:reset, Video_In_Scaler:reset]
	signal sys_reset_reset_n_ports_inv                                  : std_logic;                     -- sys_reset_reset_n:inv -> rst_controller:reset_in0

begin

	edge_detection_subsystem : component nios_system_Video_In_Subsystem_Edge_Detection_Subsystem
		port map (
			edge_detection_control_slave_address    => edge_detection_control_slave_address,                         -- edge_detection_control_slave.address
			edge_detection_control_slave_write_n    => edge_detection_control_slave_write_n,                         --                             .write_n
			edge_detection_control_slave_writedata  => edge_detection_control_slave_writedata,                       --                             .writedata
			edge_detection_control_slave_chipselect => edge_detection_control_slave_chipselect,                      --                             .chipselect
			edge_detection_control_slave_readdata   => edge_detection_control_slave_readdata,                        --                             .readdata
			sys_clk_clk                             => sys_clk_clk,                                                  --                      sys_clk.clk
			sys_reset_reset_n                       => sys_reset_reset_n,                                            --                    sys_reset.reset_n
			video_stream_sink_data                  => video_in_chroma_resampler_avalon_chroma_source_data,          --            video_stream_sink.data
			video_stream_sink_startofpacket         => video_in_chroma_resampler_avalon_chroma_source_startofpacket, --                             .startofpacket
			video_stream_sink_endofpacket           => video_in_chroma_resampler_avalon_chroma_source_endofpacket,   --                             .endofpacket
			video_stream_sink_valid                 => video_in_chroma_resampler_avalon_chroma_source_valid,         --                             .valid
			video_stream_sink_ready                 => video_in_chroma_resampler_avalon_chroma_source_ready,         --                             .ready
			video_stream_source_ready               => edge_detection_subsystem_video_stream_source_ready,           --          video_stream_source.ready
			video_stream_source_data                => edge_detection_subsystem_video_stream_source_data,            --                             .data
			video_stream_source_startofpacket       => edge_detection_subsystem_video_stream_source_startofpacket,   --                             .startofpacket
			video_stream_source_endofpacket         => edge_detection_subsystem_video_stream_source_endofpacket,     --                             .endofpacket
			video_stream_source_valid               => edge_detection_subsystem_video_stream_source_valid            --                             .valid
		);

	video_in : component nios_system_Video_In_Subsystem_Video_In
		port map (
			clk                      => sys_clk_clk,                                  --                   clk.clk
			reset                    => rst_controller_reset_out_reset,               --                 reset.reset
			stream_out_ready         => video_in_avalon_decoder_source_ready,         -- avalon_decoder_source.ready
			stream_out_startofpacket => video_in_avalon_decoder_source_startofpacket, --                      .startofpacket
			stream_out_endofpacket   => video_in_avalon_decoder_source_endofpacket,   --                      .endofpacket
			stream_out_valid         => video_in_avalon_decoder_source_valid,         --                      .valid
			stream_out_data          => video_in_avalon_decoder_source_data,          --                      .data
			TD_CLK27                 => video_in_TD_CLK27,                            --    external_interface.export
			TD_DATA                  => video_in_TD_DATA,                             --                      .export
			TD_HS                    => video_in_TD_HS,                               --                      .export
			TD_VS                    => video_in_TD_VS,                               --                      .export
			clk27_reset              => video_in_clk27_reset,                         --                      .export
			TD_RESET                 => video_in_TD_RESET,                            --                      .export
			overflow_flag            => video_in_overflow_flag                        --                      .export
		);

	video_in_csc : component nios_system_Video_In_Subsystem_Video_In_CSC
		port map (
			clk                      => sys_clk_clk,                                                --               clk.clk
			reset                    => rst_controller_reset_out_reset,                             --             reset.reset
			stream_in_startofpacket  => edge_detection_subsystem_video_stream_source_startofpacket, --   avalon_csc_sink.startofpacket
			stream_in_endofpacket    => edge_detection_subsystem_video_stream_source_endofpacket,   --                  .endofpacket
			stream_in_valid          => edge_detection_subsystem_video_stream_source_valid,         --                  .valid
			stream_in_ready          => edge_detection_subsystem_video_stream_source_ready,         --                  .ready
			stream_in_data           => edge_detection_subsystem_video_stream_source_data,          --                  .data
			stream_out_ready         => video_in_csc_avalon_csc_source_ready,                       -- avalon_csc_source.ready
			stream_out_startofpacket => video_in_csc_avalon_csc_source_startofpacket,               --                  .startofpacket
			stream_out_endofpacket   => video_in_csc_avalon_csc_source_endofpacket,                 --                  .endofpacket
			stream_out_valid         => video_in_csc_avalon_csc_source_valid,                       --                  .valid
			stream_out_data          => video_in_csc_avalon_csc_source_data                         --                  .data
		);

	video_in_chroma_resampler : component nios_system_Video_In_Subsystem_Video_In_Chroma_Resampler
		port map (
			clk                      => sys_clk_clk,                                                  --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                               --                reset.reset
			stream_in_startofpacket  => video_in_avalon_decoder_source_startofpacket,                 --   avalon_chroma_sink.startofpacket
			stream_in_endofpacket    => video_in_avalon_decoder_source_endofpacket,                   --                     .endofpacket
			stream_in_valid          => video_in_avalon_decoder_source_valid,                         --                     .valid
			stream_in_ready          => video_in_avalon_decoder_source_ready,                         --                     .ready
			stream_in_data           => video_in_avalon_decoder_source_data,                          --                     .data
			stream_out_ready         => video_in_chroma_resampler_avalon_chroma_source_ready,         -- avalon_chroma_source.ready
			stream_out_startofpacket => video_in_chroma_resampler_avalon_chroma_source_startofpacket, --                     .startofpacket
			stream_out_endofpacket   => video_in_chroma_resampler_avalon_chroma_source_endofpacket,   --                     .endofpacket
			stream_out_valid         => video_in_chroma_resampler_avalon_chroma_source_valid,         --                     .valid
			stream_out_data          => video_in_chroma_resampler_avalon_chroma_source_data           --                     .data
		);

	video_in_clipper : component nios_system_Video_In_Subsystem_Video_In_Clipper
		port map (
			clk                      => sys_clk_clk,                                            --                   clk.clk
			reset                    => rst_controller_reset_out_reset,                         --                 reset.reset
			stream_in_data           => video_in_rgb_resampler_avalon_rgb_source_data,          --   avalon_clipper_sink.data
			stream_in_startofpacket  => video_in_rgb_resampler_avalon_rgb_source_startofpacket, --                      .startofpacket
			stream_in_endofpacket    => video_in_rgb_resampler_avalon_rgb_source_endofpacket,   --                      .endofpacket
			stream_in_valid          => video_in_rgb_resampler_avalon_rgb_source_valid,         --                      .valid
			stream_in_ready          => video_in_rgb_resampler_avalon_rgb_source_ready,         --                      .ready
			stream_out_ready         => video_in_clipper_avalon_clipper_source_ready,           -- avalon_clipper_source.ready
			stream_out_data          => video_in_clipper_avalon_clipper_source_data,            --                      .data
			stream_out_startofpacket => video_in_clipper_avalon_clipper_source_startofpacket,   --                      .startofpacket
			stream_out_endofpacket   => video_in_clipper_avalon_clipper_source_endofpacket,     --                      .endofpacket
			stream_out_valid         => video_in_clipper_avalon_clipper_source_valid            --                      .valid
		);

	video_in_dma : component nios_system_Video_In_Subsystem_Video_In_DMA
		port map (
			clk                  => sys_clk_clk,                                        --                      clk.clk
			reset                => rst_controller_reset_out_reset,                     --                    reset.reset
			stream_data          => video_in_scaler_avalon_scaler_source_data,          --          avalon_dma_sink.data
			stream_startofpacket => video_in_scaler_avalon_scaler_source_startofpacket, --                         .startofpacket
			stream_endofpacket   => video_in_scaler_avalon_scaler_source_endofpacket,   --                         .endofpacket
			stream_valid         => video_in_scaler_avalon_scaler_source_valid,         --                         .valid
			stream_ready         => video_in_scaler_avalon_scaler_source_ready,         --                         .ready
			slave_address        => video_in_dma_control_slave_address,                 -- avalon_dma_control_slave.address
			slave_byteenable     => video_in_dma_control_slave_byteenable,              --                         .byteenable
			slave_read           => video_in_dma_control_slave_read,                    --                         .read
			slave_write          => video_in_dma_control_slave_write,                   --                         .write
			slave_writedata      => video_in_dma_control_slave_writedata,               --                         .writedata
			slave_readdata       => video_in_dma_control_slave_readdata,                --                         .readdata
			master_address       => video_in_dma_master_address,                        --        avalon_dma_master.address
			master_waitrequest   => video_in_dma_master_waitrequest,                    --                         .waitrequest
			master_write         => video_in_dma_master_write,                          --                         .write
			master_writedata     => video_in_dma_master_writedata                       --                         .writedata
		);

	video_in_rgb_resampler : component nios_system_Video_In_Subsystem_Video_In_RGB_Resampler
		port map (
			clk                      => sys_clk_clk,                                            --               clk.clk
			reset                    => rst_controller_reset_out_reset,                         --             reset.reset
			stream_in_startofpacket  => video_in_csc_avalon_csc_source_startofpacket,           --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => video_in_csc_avalon_csc_source_endofpacket,             --                  .endofpacket
			stream_in_valid          => video_in_csc_avalon_csc_source_valid,                   --                  .valid
			stream_in_ready          => video_in_csc_avalon_csc_source_ready,                   --                  .ready
			stream_in_data           => video_in_csc_avalon_csc_source_data,                    --                  .data
			stream_out_ready         => video_in_rgb_resampler_avalon_rgb_source_ready,         -- avalon_rgb_source.ready
			stream_out_startofpacket => video_in_rgb_resampler_avalon_rgb_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => video_in_rgb_resampler_avalon_rgb_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => video_in_rgb_resampler_avalon_rgb_source_valid,         --                  .valid
			stream_out_data          => video_in_rgb_resampler_avalon_rgb_source_data           --                  .data
		);

	video_in_scaler : component nios_system_Video_In_Subsystem_Video_In_Scaler
		port map (
			clk                      => sys_clk_clk,                                          --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                       --                reset.reset
			stream_in_startofpacket  => video_in_clipper_avalon_clipper_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => video_in_clipper_avalon_clipper_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => video_in_clipper_avalon_clipper_source_valid,         --                     .valid
			stream_in_ready          => video_in_clipper_avalon_clipper_source_ready,         --                     .ready
			stream_in_data           => video_in_clipper_avalon_clipper_source_data,          --                     .data
			stream_out_ready         => video_in_scaler_avalon_scaler_source_ready,           -- avalon_scaler_source.ready
			stream_out_startofpacket => video_in_scaler_avalon_scaler_source_startofpacket,   --                     .startofpacket
			stream_out_endofpacket   => video_in_scaler_avalon_scaler_source_endofpacket,     --                     .endofpacket
			stream_out_valid         => video_in_scaler_avalon_scaler_source_valid,           --                     .valid
			stream_out_data          => video_in_scaler_avalon_scaler_source_data             --                     .data
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_reset_reset_n_ports_inv,    -- reset_in0.reset
			clk            => sys_clk_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	sys_reset_reset_n_ports_inv <= not sys_reset_reset_n;

end architecture rtl; -- of nios_system_Video_In_Subsystem
